***************************
** fet_03v3_t_cap
***************************
* Copyright 2023 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

** library calling

.include {{model_design_path}}
.lib {{model_card_path}} {{corner}}

** Circuit Description **
* power supply
vds D_tn 0 dc={{vds_val}}
vgs G_tn 0 dc=6
vbs B_tn 0 dc={{vbs_val}}

.temp {{temp}}

* circuit
xm D_tn G_tn 0 B_tn {{device}} W = {{width}}u L = {{length}}u nf={{nf}}

.control
set filetype=ascii
set wr_singlescale
set wr_vecnames
set appendwrite

save  @m.xm.m0[vgs] @m.xm.m0[vds] @m.xm.m0[vbs] @m.xm.m0[{{cap}}]

*******************
** simulation part
*******************
DC {{main_sweep}}

* ** parameters calculation
let vgs = @m.xm.m0[vgs]
let vds = @m.xm.m0[vds]
let vbs = @m.xm.m0[vbs]
let {{cap}} = -{@m.xm.m0[{{cap}}]*1e15}

wrdata {{result_path}} vgs vds vbs {{cap}}
.endc
.end
