.SUBCKT gf180mcu_fd_io__fill1 DVDD DVSS VDD VSS
.ENDS
