.SUBCKT gf180mcu_fd_io__cor DVDD DVSS VDD VSS
C0 DVDD DVSS $[nmoscap_6p0] m=70.0 l=10e-6 w=25e-6
M1 n7 n8 VDD VDD pmos_6p0 m=1.0 w=15e-6 l=700e-9 nf=1.0 as=6.6e-12 ad=6.6e-12 
+ ps=30.88e-6 pd=30.88e-6 nrd=29.333e-3 nrs=29.333e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M2 n8 n9 VDD VDD pmos_6p0 m=1.0 w=20e-6 l=700e-9 nf=1.0 as=8.8e-12 ad=8.8e-12 
+ ps=40.88e-6 pd=40.88e-6 nrd=22e-3 nrs=22e-3 sa=440e-9 sb=440e-9 sd=0.0 
+ dtemp=0.0 par=1
M3 n5 n7 VDD VDD pmos_6p0 m=1.0 w=120e-6 l=700e-9 nf=2.0 as=52.8e-12 ad=31.2e-12 
+ ps=241.76e-6 pd=121.04e-6 nrd=2.167e-3 nrs=3.667e-3 sa=440e-9 sb=440e-9 
+ sd=520e-9 dtemp=0.0 par=1
C4 n9 VSS $[nmoscap_6p0] m=8.0 l=10e-6 w=25e-6
R5 n12 n16 $SUB=VDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R6 n11 n12 $SUB=VDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R7 n20 n11 $SUB=VDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R8 n22 n20 $SUB=VDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R9 n18 n22 $SUB=VDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R10 n21 n9 $SUB=VDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R11 n23 n21 $SUB=VDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R12 n19 n23 $SUB=VDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R13 n14 n19 $SUB=VDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R14 n13 n14 $SUB=VDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R15 n16 n13 $SUB=VDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R16 VDD n18 $SUB=VDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
M17 n8 n9 VSS VSS nmos_6p0 m=1.0 w=5e-6 l=700e-9 nf=1.0 as=2.2e-12 ad=2.2e-12 
+ ps=10.88e-6 pd=10.88e-6 nrd=88e-3 nrs=88e-3 sa=440e-9 sb=440e-9 sd=0.0 
+ dtemp=0.0 par=1
M18 VDD n5 VSS VSS nmos_6p0 m=1.0 w=4e-3 l=700e-9 nf=80.0 as=1.058e-9 ad=1.04e-9 
+ ps=4.14232e-3 pd=4.0416e-3 nrd=65e-6 nrs=66e-6 sa=440e-9 sb=440e-9 sd=520e-9 
+ dtemp=0.0 par=1
M19 n5 n7 VSS VSS nmos_6p0 m=1.0 w=30e-6 l=700e-9 nf=1.0 as=13.2e-12 ad=13.2e-12 
+ ps=60.88e-6 pd=60.88e-6 nrd=14.667e-3 nrs=14.667e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M20 n7 n8 VSS VSS nmos_6p0 m=1.0 w=30e-6 l=700e-9 nf=1.0 as=13.2e-12 ad=13.2e-12 
+ ps=60.88e-6 pd=60.88e-6 nrd=14.667e-3 nrs=14.667e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M21 n27 n28 DVDD DVDD pmos_6p0 m=1.0 w=15e-6 l=700e-9 nf=1.0 as=6.6e-12 ad=6.6e-12 
+ ps=30.88e-6 pd=30.88e-6 nrd=29.333e-3 nrs=29.333e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M22 n28 n29 DVDD DVDD pmos_6p0 m=1.0 w=20e-6 l=700e-9 nf=1.0 as=8.8e-12 ad=8.8e-12 
+ ps=40.88e-6 pd=40.88e-6 nrd=22e-3 nrs=22e-3 sa=440e-9 sb=440e-9 sd=0.0 
+ dtemp=0.0 par=1
M23 n25 n27 DVDD DVDD pmos_6p0 m=1.0 w=120e-6 l=700e-9 nf=2.0 as=52.8e-12 
+ ad=31.2e-12 ps=241.76e-6 pd=121.04e-6 nrd=2.167e-3 nrs=3.667e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
C24 n29 DVSS $[nmoscap_6p0] m=8.0 l=10e-6 w=25e-6
R25 n32 n36 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R26 n31 n32 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R27 n40 n31 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R28 n42 n40 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R29 n38 n42 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R30 n41 n29 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R31 n43 n41 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R32 n39 n43 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R33 n34 n39 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R34 n33 n34 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R35 n36 n33 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
R36 DVDD n38 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=63.855e-6 m=1.0 r=29.999e3 par=1
M37 n28 n29 DVSS DVSS nmos_6p0 m=1.0 w=5e-6 l=700e-9 nf=1.0 as=2.2e-12 ad=2.2e-12 
+ ps=10.88e-6 pd=10.88e-6 nrd=88e-3 nrs=88e-3 sa=440e-9 sb=440e-9 sd=0.0 
+ dtemp=0.0 par=1
M38 DVDD n25 DVSS DVSS nmos_6p0 m=1.0 w=4e-3 l=700e-9 nf=80.0 as=1.058e-9 ad=1.04e-9 
+ ps=4.14232e-3 pd=4.0416e-3 nrd=65e-6 nrs=66e-6 sa=440e-9 sb=440e-9 sd=520e-9 
+ dtemp=0.0 par=1
M39 n25 n27 DVSS DVSS nmos_6p0 m=1.0 w=30e-6 l=700e-9 nf=1.0 as=13.2e-12 
+ ad=13.2e-12 ps=60.88e-6 pd=60.88e-6 nrd=14.667e-3 nrs=14.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M40 n27 n28 DVSS DVSS nmos_6p0 m=1.0 w=30e-6 l=700e-9 nf=1.0 as=13.2e-12 
+ ad=13.2e-12 ps=60.88e-6 pd=60.88e-6 nrd=14.667e-3 nrs=14.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
.ENDS
