.SUBCKT gf180mcu_fd_io__fillnc DVDD DVSS VDD VSS
.ENDS
