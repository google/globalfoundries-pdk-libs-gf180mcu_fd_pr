************************************************************************
* auCdl Netlist:
* 
* Library Name:  TCG_Library
* Top Cell Name: diode_nw2ps_06v0
* View Name:     schematic
* Netlisted on:  Nov 24 09:43:35 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL vdd!

*.PIN vdd!

************************************************************************
* Library Name: TCG_Library
* Cell Name:    diode_nw2ps_06v0
* View Name:    schematic
************************************************************************

.SUBCKT diode_nw2ps_06v0 I1_0_0_0_0_R0_MINUS I1_0_1_0_0_R0_MINUS I1_0_2_0_0_R0_MINUS 
+ I1_0_3_0_0_R0_MINUS I1_1_0_0_0_R0_MINUS I1_1_1_0_0_R0_MINUS 
+ I1_1_2_0_0_R0_MINUS I1_1_3_0_0_R0_MINUS I1_2_0_0_0_R0_MINUS 
+ I1_2_1_0_0_R0_MINUS I1_2_2_0_0_R0_MINUS I1_2_3_0_0_R0_MINUS 
+ I1_3_0_0_0_R0_MINUS I1_3_1_0_0_R0_MINUS I1_3_2_0_0_R0_MINUS 
+ I1_3_3_0_0_R0_MINUS I1_default_MINUS vdd!
*.PININFO I1_0_0_0_0_R0_MINUS:I I1_0_1_0_0_R0_MINUS:I I1_0_2_0_0_R0_MINUS:I 
*.PININFO I1_0_3_0_0_R0_MINUS:I I1_1_0_0_0_R0_MINUS:I I1_1_1_0_0_R0_MINUS:I 
*.PININFO I1_1_2_0_0_R0_MINUS:I I1_1_3_0_0_R0_MINUS:I I1_2_0_0_0_R0_MINUS:I 
*.PININFO I1_2_1_0_0_R0_MINUS:I I1_2_2_0_0_R0_MINUS:I I1_2_3_0_0_R0_MINUS:I 
*.PININFO I1_3_0_0_0_R0_MINUS:I I1_3_1_0_0_R0_MINUS:I I1_3_2_0_0_R0_MINUS:I 
*.PININFO I1_3_3_0_0_R0_MINUS:I I1_default_MINUS:I vdd!:I
DI1_3_3_0_0_R0 vdd! I1_3_3_0_0_R0_MINUS diode_nw2ps_06v0 m=1 AREA=10n PJ=400u
DI1_3_2_0_0_R0 vdd! I1_3_2_0_0_R0_MINUS diode_nw2ps_06v0 m=1 AREA=1.21n PJ=224.2u
DI1_3_1_0_0_R0 vdd! I1_3_1_0_0_R0_MINUS diode_nw2ps_06v0 m=1 AREA=123p PJ=202.46u
DI1_3_0_0_0_R0 vdd! I1_3_0_0_0_R0_MINUS diode_nw2ps_06v0 m=1 AREA=86p PJ=201.72u
DI1_2_3_0_0_R0 vdd! I1_2_3_0_0_R0_MINUS diode_nw2ps_06v0 m=1 AREA=1.21n PJ=224.2u
DI1_2_2_0_0_R0 vdd! I1_2_2_0_0_R0_MINUS diode_nw2ps_06v0 m=1 AREA=146.41p PJ=48.4u
DI1_2_1_0_0_R0 vdd! I1_2_1_0_0_R0_MINUS diode_nw2ps_06v0 m=1 AREA=14.883p PJ=26.66u
DI1_2_0_0_0_R0 vdd! I1_2_0_0_0_R0_MINUS diode_nw2ps_06v0 m=1 AREA=10.406p PJ=25.92u
DI1_1_3_0_0_R0 vdd! I1_1_3_0_0_R0_MINUS diode_nw2ps_06v0 m=1 AREA=123p PJ=202.46u
DI1_1_2_0_0_R0 vdd! I1_1_2_0_0_R0_MINUS diode_nw2ps_06v0 m=1 AREA=14.883p PJ=26.66u
DI1_1_1_0_0_R0 vdd! I1_1_1_0_0_R0_MINUS diode_nw2ps_06v0 m=1 AREA=1.5129p PJ=4.92u
DI1_1_0_0_0_R0 vdd! I1_1_0_0_0_R0_MINUS diode_nw2ps_06v0 m=1 AREA=1.0578p PJ=4.18u
DI1_0_3_0_0_R0 vdd! I1_0_3_0_0_R0_MINUS diode_nw2ps_06v0 m=1 AREA=86p PJ=201.72u
DI1_0_2_0_0_R0 vdd! I1_0_2_0_0_R0_MINUS diode_nw2ps_06v0 m=1 AREA=10.406p PJ=25.92u
DI1_0_1_0_0_R0 vdd! I1_0_1_0_0_R0_MINUS diode_nw2ps_06v0 m=1 AREA=1.0578p PJ=4.18u
DI1_0_0_0_0_R0 vdd! I1_0_0_0_0_R0_MINUS diode_nw2ps_06v0 m=1 AREA=739.6f PJ=3.44u
DI1_default vdd! I1_default_MINUS diode_nw2ps_06v0 m=1 AREA=1p PJ=4u
.ENDS

