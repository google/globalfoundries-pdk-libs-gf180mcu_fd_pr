*Xyce Common Source Circuit
** library calling



*****************
** main netlist
*****************

Vcp c 0 dc 6
Ib 0 b 9u

xq1 c b 0 0 vnpn_10x10


*****************
** Analysis
*****************
.DC Vcp 0 6 0.1 Ib 1u 9u 2u
.STEP TEMP 25 -60 200
.print DC FORMAT=CSV file=result.csv {-I(Vcp)}

.include "../../design.xyce"
.lib "../../sm141064.xyce" bjt_typical

.end
