***************************
** nfet_03v3_t_id
***************************
* Copyright 2022 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
Vds D_tn 0 dc -6.6
Vgs G_tn 0 -6

.temp 25
.options tnom=25

xmn1 D_tn G_tn 0 0 pfet_06v0_dss W = 5u L = 1.0u ad=1.2u pd=10.48u as=1.2u ps=10.48u

**** begin architecture code


.control
set filetype=ascii

dc Vds 0 -6.6 -0.05 Vgs -1 -6 -1
print i(Vds)
wrdata mos_iv_regr/pfet_06v0_dss_iv/simulated_Id/T25_simulated_W5_L1.0.csv i(Vds)
.endc



** library calling

.include "../../../design.ngspice"
.lib "../../../sm141064.ngspice" typical


**** end architecture code


.end