************************************************************************
* auCdl Netlist:
* 
* Library Name:  TCG_Library
* Top Cell Name: vpnp_10x10
* View Name:     schematic
* Netlisted on:  Nov 24 10:36:53 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: TCG_Library
* Cell Name:    vpnp_10x10
* View Name:    schematic
************************************************************************

.SUBCKT vpnp_10x10 I1_default_B I1_default_C I1_default_E
*.PININFO I1_default_B:I I1_default_C:I I1_default_E:I
QI1_default I1_default_C I1_default_B I1_default_E vpnp_10x10 m=1
.ENDS

