*Xyce Common Source Circuit
** library calling


*****************
** main netlist
*****************
Vn n 0 dc 1


dn1 n 0 {{device}} AREA={{area}}p
* PJ=40u


*****************
** Analysis
*****************
.DC Vn -40.41 1.41 0.41
.STEP TEMP {{temp}} -60 200
.print DC FORMAT=CSV file=diode_regr/{{device}}/simulated_iv/simulated_A{{area}}_P{{pj}}_t{{temp}}_{{corner}}.csv {abs(I(dn1))}

* .print DC FORMAT=CSV file=result.csv {N(dn1:is)}




.include "../../../design.xyce"
.lib "../../../sm141064.xyce" diode_{{corner}}

.end
