******************
** MIMCAP NETLISTS
******************
* Copyright 2023 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

*****************
** main netlist
*****************
.param volt = -3.0

V1 in 0 dc {volt} ac 1
R1 in out 1G
xcn out 0 {{device}} c_length={{length}}u c_width={{width}}u l={{length}}u w={{width}}u

.meas AC freq when Vdb(out)=-3 PRECISION=15

*****************
** Analysis
*****************

.ac dec 10 1 10G
.step volt {{voltage}}

.include {{model_design_path}}
.lib {{model_card_path}} {{corner}}

.end
