****************
** cap_mos_cv **
****************
* Copyright 2023 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
.options noacct

.ic v(cc)=0.0

.temp {{temp}}

Vinp inp 0 dc={{supp_val}}
R1 inp cc {{res_val}}k
xcn cc 0 {{device}} c_length={{length}}u c_width={{width}}u

.control
    ** unset askquit
    tran 50ps {{sim_run_time}}ps uic
    let q_t = integ(-i(vinp))
    wrdata {{result_path_pos}} v(cc) q_t

    alter vinp dc=-{{supp_val}}
    tran 50ps {{sim_run_time}}ps uic
    let q_t = integ(-i(vinp))
    wrdata {{result_path_neg}} v(cc) q_t
.endc

** library calling

.include "../../../design.ngspice"
.lib "../../../sm141064.ngspice" {{corner}}
.end
