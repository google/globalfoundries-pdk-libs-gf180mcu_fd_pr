*Xyce Common Source Circuit
** library calling


*****************
** main netlist
*****************
Vds D_tn 0 dc 0.05
Vgs G_tn 0 dc 3.3
Vbs S_tn 0 dc 0

xmn1 D_tn G_tn 0 S_tn nmos_3p3 W=10u L=10u ad=2.4u pd=20.48u as=2.4u ps=20.48u


*****************
** Analysis
*****************
.dc Vgs 0 3.3 0.05 Vbs 0 -3.3 -0.825
.STEP TEMP -40 -60 200
.print DC FORMAT=CSV file=result.csv {-I(Vds)}

.include "../../../../design.xyce"
.lib "../../../../sm141064.xyce" typical

.end
