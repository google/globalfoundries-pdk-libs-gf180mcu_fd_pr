.SUBCKT gf180mcu_fd_io__bi_t A CS DVDD DVSS IE OE PAD PD PDRV0 PDRV1 PU SL VDD VSS Y
C0 DVDD DVSS $[nmoscap_6p0] m=4.0 l=3e-6 w=3e-6
C1 DVDD DVSS $[nmoscap_6p0] m=10.0 l=1.5e-6 w=5e-6
M2 n67 n75 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 ad=1.32e-12 
+ ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M3 n37 n67 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 ad=1.32e-12 
+ ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M4 n72 OE VSS VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 ad=1.32e-12 
+ ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M5 n75 A n72 VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M6 n67 n75 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 ad=2.64e-12 
+ ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M7 n37 n67 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 ad=2.64e-12 
+ ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M8 n75 OE VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 ad=1.32e-12 
+ ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M9 n75 A VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 ad=1.32e-12 
+ ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M10 PAD n43 DVDD DVDD pmos_6p0_sab m=1.0 w=80e-6 l=700e-9 nf=2.0 s_sab=280e-9 
+ d_sab=2.78e-6 par=1 dtemp=0.0
M11 PAD n55 DVSS DVSS nmos_6p0_sab m=1.0 w=38e-6 l=1.15e-6 nf=1.0 s_sab=280e-9 
+ d_sab=3.78e-6 par=1 dtemp=0.0
M12 PAD n52 DVSS DVSS nmos_6p0_sab m=1.0 w=38e-6 l=1.15e-6 nf=1.0 s_sab=280e-9 
+ d_sab=3.78e-6 par=1 dtemp=0.0
M13 PAD n48 DVDD DVDD pmos_6p0_sab m=1.0 w=40e-6 l=700e-9 nf=1.0 s_sab=280e-9 
+ d_sab=2.78e-6 par=1 dtemp=0.0
M14 PAD n42 DVDD DVDD pmos_6p0_sab m=1.0 w=80e-6 l=700e-9 nf=2.0 s_sab=280e-9 
+ d_sab=2.78e-6 par=1 dtemp=0.0
M15 PAD n56 DVSS DVSS nmos_6p0_sab m=1.0 w=38e-6 l=1.15e-6 nf=1.0 s_sab=280e-9 
+ d_sab=3.78e-6 par=1 dtemp=0.0
M16 PAD n51 DVSS DVSS nmos_6p0_sab m=1.0 w=38e-6 l=1.15e-6 nf=1.0 s_sab=280e-9 
+ d_sab=3.78e-6 par=1 dtemp=0.0
M17 PAD n47 DVDD DVDD pmos_6p0_sab m=1.0 w=40e-6 l=700e-9 nf=1.0 s_sab=280e-9 
+ d_sab=2.78e-6 par=1 dtemp=0.0
M18 PAD n44 DVDD DVDD pmos_6p0_sab m=1.0 w=80e-6 l=700e-9 nf=2.0 s_sab=280e-9 
+ d_sab=2.78e-6 par=1 dtemp=0.0
M19 PAD n54 DVSS DVSS nmos_6p0_sab m=1.0 w=38e-6 l=1.15e-6 nf=1.0 s_sab=280e-9 
+ d_sab=3.78e-6 par=1 dtemp=0.0
M20 PAD n53 DVSS DVSS nmos_6p0_sab m=1.0 w=38e-6 l=1.15e-6 nf=1.0 s_sab=280e-9 
+ d_sab=3.78e-6 par=1 dtemp=0.0
M21 PAD n49 DVDD DVDD pmos_6p0_sab m=1.0 w=40e-6 l=700e-9 nf=1.0 s_sab=280e-9 
+ d_sab=2.78e-6 par=1 dtemp=0.0
M22 PAD n45 DVDD DVDD pmos_6p0_sab m=1.0 w=80e-6 l=700e-9 nf=2.0 s_sab=280e-9 
+ d_sab=2.78e-6 par=1 dtemp=0.0
M23 PAD n57 DVSS DVSS nmos_6p0_sab m=1.0 w=38e-6 l=1.15e-6 nf=1.0 s_sab=280e-9 
+ d_sab=3.78e-6 par=1 dtemp=0.0
M24 PAD n50 DVSS DVSS nmos_6p0_sab m=1.0 w=38e-6 l=1.15e-6 nf=1.0 s_sab=280e-9 
+ d_sab=3.78e-6 par=1 dtemp=0.0
M25 PAD n46 DVDD DVDD pmos_6p0_sab m=1.0 w=40e-6 l=700e-9 nf=1.0 s_sab=280e-9 
+ d_sab=2.78e-6 par=1 dtemp=0.0
M26 n58 n41 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 ad=780e-15 
+ ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9 
+ sd=520e-9 dtemp=0.0 par=1
M27 n175 SL VSS VSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M28 n41 n175 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M29 n58 n41 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M30 n175 SL VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M31 n41 n175 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
D32 A VDD pn_6p0 m=1.0 AREA=1e-12 PJ=4e-6
D33 SL VDD pn_6p0 m=1.0 AREA=1e-12 PJ=4e-6
D34 VSS PDRV0 pn_6p0 m=1.0 AREA=230.4e-15 PJ=1.92e-6
D35 VSS OE pn_6p0 m=1.0 AREA=230.4e-15 PJ=1.92e-6
M36 n188 PDRV0 VSS VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M37 n179 OE n188 VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M38 n39 n36 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M39 n36 n179 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M40 n179 PDRV0 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M41 n179 OE VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M42 n39 n36 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M43 n36 n179 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
D44 VSS PDRV1 pn_6p0 m=1.0 AREA=230.4e-15 PJ=1.92e-6
D45 VSS OE pn_6p0 m=1.0 AREA=230.4e-15 PJ=1.92e-6
M46 n198 PDRV1 VSS VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M47 n189 OE n198 VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M48 n35 n33 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M49 n33 n189 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M50 n189 PDRV1 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M51 n189 OE VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M52 n35 n33 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M53 n33 n189 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
D54 VSS VDD pn_6p0 m=1.0 AREA=230.4e-15 PJ=1.92e-6
D55 VSS OE pn_6p0 m=1.0 AREA=230.4e-15 PJ=1.92e-6
M56 n208 VDD VSS VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M57 n199 OE n208 VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M58 n32 n31 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M59 n31 n199 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M60 n199 VDD VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M61 n199 OE VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M62 n32 n31 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M63 n31 n199 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M64 n46 n58 n45 DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M65 n45 DVDD n46 DVSS nmos_6p0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15 
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M66 n50 n209 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M67 n57 n209 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M68 n46 n214 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M69 n214 n37 DVSS DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M70 n214 n39 DVSS DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M71 n209 n36 n214 DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M72 n50 n41 n57 DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M73 n209 n36 DVDD DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M74 n46 n214 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M75 n57 n209 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M76 n50 DVSS n57 DVDD pmos_6p0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15 
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M77 n209 n37 DVDD DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M78 n214 n39 n209 DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M79 n45 n214 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M80 n47 n58 n42 DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M81 n42 DVDD n47 DVSS nmos_6p0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15 
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M82 n51 n222 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M83 n56 n222 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M84 n47 n227 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M85 n227 n37 DVSS DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M86 n227 n35 DVSS DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M87 n222 n33 n227 DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M88 n51 n41 n56 DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M89 n222 n33 DVDD DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M90 n47 n227 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M91 n56 n222 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M92 n51 DVSS n56 DVDD pmos_6p0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15 
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M93 n222 n37 DVDD DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M94 n227 n35 n222 DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M95 n42 n227 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M96 n48 n58 n43 DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M97 n43 DVDD n48 DVSS nmos_6p0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15 
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M98 n52 n235 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M99 n55 n235 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M100 n48 n240 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M101 n240 n37 DVSS DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M102 n240 n35 DVSS DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M103 n235 n33 n240 DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M104 n52 n41 n55 DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M105 n235 n33 DVDD DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M106 n48 n240 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M107 n55 n235 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M108 n52 DVSS n55 DVDD pmos_6p0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15 
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M109 n235 n37 DVDD DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M110 n240 n35 n235 DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M111 n43 n240 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M112 n49 n58 n44 DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M113 n44 DVDD n49 DVSS nmos_6p0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15 
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M114 n53 n248 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M115 n54 n248 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M116 n49 n253 DVSS DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M117 n253 n37 DVSS DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M118 n253 n32 DVSS DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M119 n248 n31 n253 DVSS nmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M120 n53 n41 n54 DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M121 n248 n31 DVDD DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M122 n49 n253 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M123 n54 n248 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M124 n53 DVSS n54 DVDD pmos_6p0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15 
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M125 n248 n37 DVDD DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M126 n253 n32 n248 DVDD pmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M127 n44 n253 DVDD DVDD pmos_6p0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M128 n273 n262 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M129 n286 IE VSS VSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M130 n262 n286 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M131 n273 n262 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M132 n286 IE VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M133 n262 n286 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M134 n279 n263 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M135 n294 CS VSS VSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M136 n263 n294 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M137 n279 n263 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M138 n294 CS VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M139 n263 n294 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M140 n277 n265 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M141 n302 n266 VSS VSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M142 n265 n302 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M143 n277 n265 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M144 n302 n266 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M145 n265 n302 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M146 n281 n268 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M147 n310 n264 VSS VSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M148 n268 n310 DVSS DVSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M149 n281 n268 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M150 n310 n264 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M151 n268 n310 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
D152 PD VDD pn_6p0 m=1.0 AREA=1e-12 PJ=4e-6
D153 IE VDD pn_6p0 m=1.0 AREA=1e-12 PJ=4e-6
D154 CS VDD pn_6p0 m=1.0 AREA=1e-12 PJ=4e-6
D155 PU VDD pn_6p0 m=1.0 AREA=1e-12 PJ=4e-6
M156 n318 n263 DVDD DVDD pmos_6p0 m=1.0 w=8e-6 l=700e-9 nf=1.0 as=3.52e-12 
+ ad=3.52e-12 ps=16.88e-6 pd=16.88e-6 nrd=55e-3 nrs=55e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M157 DVDD n263 n319 DVDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M158 n320 n20 DVDD DVDD pmos_6p0 m=1.0 w=3.8e-6 l=700e-9 nf=1.0 as=1.672e-12 
+ ad=1.672e-12 ps=8.48e-6 pd=8.48e-6 nrd=115.789e-3 nrs=115.789e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M159 DVSS n319 n320 DVDD pmos_6p0 m=1.0 w=3.8e-6 l=700e-9 nf=1.0 as=1.672e-12 
+ ad=1.672e-12 ps=8.48e-6 pd=8.48e-6 nrd=115.789e-3 nrs=115.789e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M160 n280 n262 DVDD DVDD pmos_6p0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M161 n280 n318 n315 DVDD pmos_6p0 m=1.0 w=2e-6 l=700e-9 nf=1.0 as=880e-15 
+ ad=880e-15 ps=4.88e-6 pd=4.88e-6 nrd=220e-3 nrs=220e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M162 n280 n318 n319 DVDD pmos_6p0 m=1.0 w=2e-6 l=700e-9 nf=1.0 as=880e-15 
+ ad=880e-15 ps=4.88e-6 pd=4.88e-6 nrd=220e-3 nrs=220e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M163 n280 n20 n320 DVDD pmos_6p0 m=1.0 w=4.3e-6 l=700e-9 nf=1.0 as=1.892e-12 
+ ad=1.892e-12 ps=9.48e-6 pd=9.48e-6 nrd=102.326e-3 nrs=102.326e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M164 n325 n262 DVSS DVSS nmos_6p0 m=1.0 w=16e-6 l=700e-9 nf=1.0 as=7.04e-12 
+ ad=7.04e-12 ps=32.88e-6 pd=32.88e-6 nrd=27.5e-3 nrs=27.5e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M165 n317 n20 n325 DVSS nmos_6p0 m=1.0 w=10.6e-6 l=700e-9 nf=1.0 as=4.664e-12 
+ ad=4.664e-12 ps=22.08e-6 pd=22.08e-6 nrd=41.509e-3 nrs=41.509e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M166 n280 n20 n317 DVSS nmos_6p0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M167 n318 n263 DVSS DVSS nmos_6p0 m=1.0 w=4e-6 l=700e-9 nf=1.0 as=1.76e-12 
+ ad=1.76e-12 ps=8.88e-6 pd=8.88e-6 nrd=110e-3 nrs=110e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M168 n280 n263 n315 DVSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M169 n280 n263 n319 DVSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M170 DVDD n315 n317 DVSS nmos_6p0 m=1.0 w=1.3e-6 l=700e-9 nf=1.0 as=572e-15 
+ ad=572e-15 ps=3.48e-6 pd=3.48e-6 nrd=338.462e-3 nrs=338.462e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M171 DVSS n318 n315 DVSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M172 n333 n280 DVDD DVDD pmos_6p0 m=1.0 w=2e-6 l=700e-9 nf=1.0 as=880e-15 
+ ad=880e-15 ps=4.88e-6 pd=4.88e-6 nrd=220e-3 nrs=220e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M173 n330 n333 VDD VDD pmos_6p0 m=1.0 w=10e-6 l=700e-9 nf=1.0 as=4.4e-12 
+ ad=4.4e-12 ps=20.88e-6 pd=20.88e-6 nrd=44e-3 nrs=44e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M174 Y n330 VDD VDD pmos_6p0 m=1.0 w=21e-6 l=700e-9 nf=1.0 as=9.24e-12 
+ ad=9.24e-12 ps=42.88e-6 pd=42.88e-6 nrd=20.952e-3 nrs=20.952e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M175 n333 n280 DVSS DVSS nmos_6p0 m=1.0 w=8e-6 l=700e-9 nf=1.0 as=3.52e-12 
+ ad=3.52e-12 ps=16.88e-6 pd=16.88e-6 nrd=55e-3 nrs=55e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M176 Y n330 VSS VSS nmos_6p0 m=1.0 w=9e-6 l=700e-9 nf=1.0 as=3.96e-12 
+ ad=3.96e-12 ps=18.88e-6 pd=18.88e-6 nrd=48.889e-3 nrs=48.889e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M177 n330 n333 VSS VSS nmos_6p0 m=1.0 w=2.5e-6 l=700e-9 nf=1.0 as=1.1e-12 
+ ad=1.1e-12 ps=5.88e-6 pd=5.88e-6 nrd=176e-3 nrs=176e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M178 n266 n340 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M179 n266 PU VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M180 n341 PU VSS VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M181 n266 n340 n341 VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M182 n264 PD VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M183 n264 n340 VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M184 n347 n340 VSS VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M185 n264 PD n347 VSS nmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M186 n353 n359 n340 VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M187 PU PD n340 VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M188 n359 PD VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M189 n353 PU VDD VDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M190 n353 PD n340 VSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M191 PU n359 n340 VSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M192 n359 PD VSS VSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M193 n353 PU VSS VSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
R194 n20 n362 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=23e-6 m=1.0 r=9.94533e3 par=1
R195 n362 n361 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
R196 n361 n360 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
R197 n360 n363 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
R198 n363 n368 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
R199 n368 n367 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
R200 n367 n364 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
R201 n364 n365 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
M202 n365 n281 DVSS DVSS nmos_6p0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M203 n365 n265 DVDD DVDD pmos_6p0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
D204 DVSS n20 np_6p0 m=2.0 AREA=20e-12 PJ=42e-6
D205 n20 DVDD pn_6p0 m=2.0 AREA=20e-12 PJ=42e-6
R206 PAD n20 $SUB=DVDD $[ppolyf_u] $W=2.5e-6 $L=2.8e-6 m=1.0 r=432.59 par=1
R207 PAD n20 $SUB=DVDD $[ppolyf_u] $W=2.5e-6 $L=2.8e-6 m=1.0 r=449.157 par=1
R208 PAD n20 $SUB=DVDD $[ppolyf_u] $W=2.5e-6 $L=2.8e-6 m=1.0 r=432.59 par=1
R209 PAD n20 $SUB=DVDD $[ppolyf_u] $W=2.5e-6 $L=2.8e-6 m=1.0 r=449.157 par=1
.ENDS
