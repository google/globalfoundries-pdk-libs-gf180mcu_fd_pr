************************************************************************
* auCdl Netlist:
* 
* Library Name:  TCG_Library
* Top Cell Name: rm3
* View Name:     schematic
* Netlisted on:  Nov 24 10:17:35 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: TCG_Library
* Cell Name:    rm3
* View Name:    schematic
************************************************************************

.SUBCKT rm3
*.PININFO
RI1_2_2_R0 net1 net2 rm3 W=50u L=50u m=1 r=90m dtemp=0
RI1_2_1_R0 net3 net4 rm3 W=50u L=13.5u m=1 r=24.3m dtemp=0
RI1_2_0_R0 net5 net6 rm3 W=50u L=280n m=1 r=504u dtemp=0
RI1_1_2_R0 net7 net8 rm3 W=13.5u L=50u m=1 r=333.333m dtemp=0
RI1_1_1_R0 net9 net10 rm3 W=13.5u L=13.5u m=1 r=90m dtemp=0
RI1_1_0_R0 net11 net12 rm3 W=13.5u L=280n m=1 r=1.86667m dtemp=0
RI1_0_2_R0 net13 net14 rm3 W=280n L=50u m=1 r=16.0714 dtemp=0
RI1_0_1_R0 net15 net16 rm3 W=280n L=13.5u m=1 r=4.33929 dtemp=0
RI1_0_0_R0 net17 net18 rm3 W=280n L=280n m=1 r=90m dtemp=0
RI1_default net19 net20 rm3 W=280.00n L=280.00n m=1 r=90.00m dtemp=0
.ENDS

