******************
** MIMCAP NETLISTS
******************
* Copyright 2023 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

Ich 0 p dc 1n

.STEP TEMP LIST {{temp}}
      
xcn p 0 {{device}} c_length={{length}}u c_width={{width}}u

.ic v(p)=0.0
.tran 1ns 10ns

.meas tran cj FIND par('(1.0e-9  * time / v(p))*1.0e15') AT=10ns


** library calling

.include {{model_design_path}}
.lib {{model_card_path}} {{corner}}

.end
