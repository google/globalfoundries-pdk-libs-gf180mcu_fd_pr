*Xyce Common Source Circuit
** library calling



*****************
** main netlist
*****************

Vcp c 0 dc -6
Ib f b -9u
Vbp f 0 dc 0
xq1 c b 0 {{device}}


*****************
** Analysis
*****************
.DC Vcp 0 -3 -0.1 Ib -1u -9u -2u
.STEP TEMP {{temp}} -60 200
.print DC FORMAT=CSV file=bjt_iv_reg/pnp/simulated/t{{temp}}_simulated_{{device}}.csv {I(Vcp)} i(Vbp) v(c)

.include "../../../../../../design.xyce"
.lib "../../../../../../sm141064.xyce" bjt_typical

.end
