*******************
** BJT-beta netlist
*******************
* Copyright 2023 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

Vcp c 0 dc=3
Vbp b 0 dc=1.2

.temp {{temp}}

xq {{terminals}} {{device}}

*****************
** Analysis
*****************
.control
set filetype=ascii
set wr_singlescale
set wr_vecnames

dc {{sweep}}

let vcp = v(c)
let vbp = v(b)
let ic = abs(-i(Vcp))
let ib = abs(-i(Vbp))

wrdata {{result_path}} vcp vbp  ic ib
.endc

** library calling

.include "../../../design.ngspice"
.lib "../../../sm141064.ngspice" {{corner}}

**** end architecture code

.end
