***************************
** nfet_06v0_t_id
***************************
* Copyright 2022 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
* power supply
Vds D_tn 0 dc=0.05
Vgs G_tn 0 dc=6
Vbs S_tn 0 dc=0

.temp {{temp}}
.options tnom={{temp}}

xmn1 D_tn G_tn 0 S_tn nfet_06v0 W = {{width}}u L = {{length}}u

**** begin architecture code


.control
set filetype=ascii

dc Vgs 0 6 0.05 Vbs 0 -3 -0.75
print -i(Vds)
wrdata nfet_06v0_iv/simulated_Id/{{i}}_simulated_W{{width}}_L{{length}}.csv -i(Vds)
.endc



** library calling

.include "../../../design.ngspice"
.lib "../../../sm141064.ngspice" typical

**** end architecture code


.end
