*Xyce Common Source Circuit
** library calling



*****************
** main netlist
*****************
Vds D_tn 0 dc 3.3
Vgs G_tn 0 dc 3.3


xmn1 D_tn G_tn 0 0 nfet_03v3 W=10u L=10u ad=2.4u pd=20.48u as=2.4u ps=20.48u



*****************
** Analysis
*****************
.DC Vds 0 3.3 0.05 Vgs 0.8 3.3 0.5
.STEP TEMP -40 -40 -40
.print DC FORMAT=CSV file=result.csv {1/N(xmn1:m0:gds)}

.include "../../design.xyce"
.lib "../../sm141064.xyce" typical

.end