.SUBCKT gf180mcu_fd_io__brk2 VSS
.ENDS
