***************************
** nfet_03v3_cv
***************************
* Copyright 2022 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
** library calling

.include "../../../design.ngspice"
.lib "../../../sm141064.ngspice" typical


** Circuit Description **
* power supply
vds D_tn 0 dc=3.3
vgs G_tn 0 dc=3.3
vs S_tn 0 dc=0

.temp 25
.options tnom=25

*l_diff_min = 0.24
* ad = int((nf+1)/2) * width/nf * 0.24       = 24u                         
* pd = (int((nf+1)/2) * width/nf + 0.24)*2   = 200.48u                 

* circuit
xmn D_tn G_tn S_tn S_tn nfet_06v0_dss W = {{width}}u L = {{length}}u nf={{nf}} ad= 24u pd=200.48u as=24u ps=200.48u

.control
set filetype=ascii

let vds_min  = 0
let vds_step = 0.1
let vds_max  = 3.3

compose  vgs_vector   start=0          stop=3.3          step=1

set appendwrite

foreach t 25

    let vgs_counter = 0
    while vgs_counter < length(vgs_vector)
        option TEMP=25
        alter vgs = vgs_vector[vgs_counter]

        save  @m.xmn.m0[vds] @m.xmn.m0[vgs] @m.xmn.m0[id] @m.xmn.m0[cgs]
        *******************
        ** simulation part
        *******************
        DC vds $&vds_min $&vds_max $&vds_step
    
        * ** parameters calculation
	
	print @m.xmn.m0[cgs]
        
        wrdata mos_cv_regr/nfet_06v0_dss/simulated_Cgs/simulated_W{{width}}_L{{length}}.csv -{@m.xmn.m0[cgs]*1e15} 
        
        reset
        let vgs_counter = vgs_counter + 1
    end
end
.endc
.end
