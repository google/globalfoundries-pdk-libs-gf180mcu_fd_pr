***************************
** nfet_06v0_nvt_t_id
***************************
* Copyright 2022 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
Vds D_tn 0 dc 6.6
Vgs G_tn 0 6

.temp 125
.options tnom=125

xmn1 D_tn G_tn 0 0 nfet_06v0_nvt W = 10u L = 10.0u ad=2.4u pd=20.48u as=2.4u ps=20.48u

**** begin architecture code


.control
set filetype=ascii

dc Vds 0 6.6 0.05 Vgs 0.25 6 1.15
print -i(Vds)
wrdata mos_iv_regr/nfet_06v0_nvt_iv/simulated_Id/T125_simulated_W10_L10.0.csv -i(Vds)
.endc



** library calling

.include "../../../design.ngspice"
.lib "../../../sm141064.ngspice" typical

**** end architecture code


.end