************************************************************************
* auCdl Netlist:
* 
* Library Name:  TCG_Library
* Top Cell Name: dnwpw_6p0
* View Name:     schematic
* Netlisted on:  Nov 24 09:07:04 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL vdd!

*.PIN vdd!

************************************************************************
* Library Name: TCG_Library
* Cell Name:    dnwpw_6p0
* View Name:    schematic
************************************************************************

.SUBCKT dnwpw_6p0 I1_0_0_0_0_R0_POS I1_0_1_0_0_R0_POS I1_0_2_0_0_R0_POS 
+ I1_1_0_0_0_R0_POS I1_1_1_0_0_R0_POS I1_1_2_0_0_R0_POS I1_2_0_0_0_R0_POS 
+ I1_2_1_0_0_R0_POS I1_2_2_0_0_R0_POS I1_default_POS vdd!
*.PININFO I1_0_0_0_0_R0_POS:I I1_0_1_0_0_R0_POS:I I1_0_2_0_0_R0_POS:I 
*.PININFO I1_1_0_0_0_R0_POS:I I1_1_1_0_0_R0_POS:I I1_1_2_0_0_R0_POS:I 
*.PININFO I1_2_0_0_0_R0_POS:I I1_2_1_0_0_R0_POS:I I1_2_2_0_0_R0_POS:I 
*.PININFO I1_default_POS:I vdd!:I
DI1_2_2_0_0_R0 I1_2_2_0_0_R0_POS vdd! dnwpw_6p0 10n 400e-6 m=1
DI1_2_1_0_0_R0 I1_2_1_0_0_R0_POS vdd! dnwpw_6p0 1.023n 220.46e-6 m=1
DI1_2_0_0_0_R0 I1_2_0_0_0_R0_POS vdd! dnwpw_6p0 74p 201.48e-6 m=1
DI1_1_2_0_0_R0 I1_1_2_0_0_R0_POS vdd! dnwpw_6p0 1.023n 220.46e-6 m=1
DI1_1_1_0_0_R0 I1_1_1_0_0_R0_POS vdd! dnwpw_6p0 104.653p 40.92e-6 m=1
DI1_1_0_0_0_R0 I1_1_0_0_0_R0_POS vdd! dnwpw_6p0 7.5702p 21.94e-6 m=1
DI1_0_2_0_0_R0 I1_0_2_0_0_R0_POS vdd! dnwpw_6p0 74p 201.48e-6 m=1
DI1_0_1_0_0_R0 I1_0_1_0_0_R0_POS vdd! dnwpw_6p0 7.5702p 21.94e-6 m=1
DI1_0_0_0_0_R0 I1_0_0_0_0_R0_POS vdd! dnwpw_6p0 595.7f 3.09e-6 m=1
DI1_default I1_default_POS vdd! dnwpw_6p0 100e-12 40e-6 m=1
.ENDS

