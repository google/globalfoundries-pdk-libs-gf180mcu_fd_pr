************************************************************************
* auCdl Netlist:
* 
* Library Name:  TCG_Library
* Top Cell Name: dnwps_3p3
* View Name:     schematic
* Netlisted on:  Nov 24 09:04:18 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL gnd!

*.PIN gnd!

************************************************************************
* Library Name: TCG_Library
* Cell Name:    dnwps_3p3
* View Name:    schematic
************************************************************************

.SUBCKT dnwps_3p3 I1_0_0_0_0_R0_NEG I1_0_1_0_0_R0_NEG I1_0_2_0_0_R0_NEG 
+ I1_1_0_0_0_R0_NEG I1_1_1_0_0_R0_NEG I1_1_2_0_0_R0_NEG I1_2_0_0_0_R0_NEG 
+ I1_2_1_0_0_R0_NEG I1_2_2_0_0_R0_NEG I1_default_NEG gnd!
*.PININFO I1_0_0_0_0_R0_NEG:I I1_0_1_0_0_R0_NEG:I I1_0_2_0_0_R0_NEG:I 
*.PININFO I1_1_0_0_0_R0_NEG:I I1_1_1_0_0_R0_NEG:I I1_1_2_0_0_R0_NEG:I 
*.PININFO I1_2_0_0_0_R0_NEG:I I1_2_1_0_0_R0_NEG:I I1_2_2_0_0_R0_NEG:I 
*.PININFO I1_default_NEG:I gnd!:I
DI1_2_2_0_0_R0 gnd! I1_2_2_0_0_R0_NEG dnwps_3p3 10n 400e-6 m=1
DI1_2_1_0_0_R0 gnd! I1_2_1_0_0_R0_NEG dnwps_3p3 1.034n 220.68e-6 m=1
DI1_2_0_0_0_R0 gnd! I1_2_0_0_0_R0_NEG dnwps_3p3 170p 203.4e-6 m=1
DI1_1_2_0_0_R0 gnd! I1_1_2_0_0_R0_NEG dnwps_3p3 1.034n 220.68e-6 m=1
DI1_1_1_0_0_R0 gnd! I1_1_1_0_0_R0_NEG dnwps_3p3 106.916p 41.36e-6 m=1
DI1_1_0_0_0_R0 gnd! I1_1_0_0_0_R0_NEG dnwps_3p3 17.578p 24.08e-6 m=1
DI1_0_2_0_0_R0 gnd! I1_0_2_0_0_R0_NEG dnwps_3p3 170p 203.4e-6 m=1
DI1_0_1_0_0_R0 gnd! I1_0_1_0_0_R0_NEG dnwps_3p3 17.578p 24.08e-6 m=1
DI1_0_0_0_0_R0 gnd! I1_0_0_0_0_R0_NEG dnwps_3p3 3.1535p 7.11e-6 m=1
DI1_default gnd! I1_default_NEG dnwps_3p3 100e-12 40e-6 m=1
.ENDS

