* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* Sources
Vdd VDD 0 dc 5
Vin1 I1 0 dc pulse(0 5 200p 1p 1p 200p 400p)
Vin2 I2 0 dc pulse(0 5 400p 1p 1p 400p 800p)
Vin3 I3 0 dc pulse(0 5 800p 1p 1p 800p 1600p)

* Main circuit
X1 I1 I2 I3 ZN VDD VDD 0 0 gf180mcu_fd_sc_mcu7t5v0__or3_1

* Temperature set
.temp 25
.options tnom=25

* Analyses
.control
tran 1p 1600p
meas tran o0 FIND V(ZN) AT=200p
meas tran o1 FIND V(ZN) AT=400p
meas tran o2 FIND V(ZN) AT=600p
meas tran o3 FIND V(ZN) AT=800p
meas tran o4 FIND V(ZN) AT=1000p
meas tran o5 FIND V(ZN) AT=1200p
meas tran o6 FIND V(ZN) AT=1400p
meas tran o7 FIND V(ZN) AT=1600p

wrdata or3/or3_simulated.csv {o0} {o1} {o2} {o3} {o4} {o5} {o6} {o7}
.endc

* Libraries calling
.include "../../../../design.xyce"
.lib "../../../../sm141064.xyce" typical

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
M_i_2 VSS A1 Z_neg VPW nmos_6p0 W=4e-07 L=6e-07
M_i_3 Z_neg A2 VSS VPW nmos_6p0 W=4e-07 L=6e-07
M_i_4 VSS A3 Z_neg VPW nmos_6p0 W=4e-07 L=6e-07
M_i_0 Z Z_neg VSS VPW nmos_6p0 W=8.2e-07 L=6e-07
M_i_5 net_0 A1 Z_neg VNW pmos_6p0 W=5.6e-07 L=5e-07
M_i_6 net_1 A2 net_0 VNW pmos_6p0 W=5.6e-07 L=5e-07
M_i_7 VDD A3 net_1 VNW pmos_6p0 W=5.6e-07 L=5e-07
M_i_1 Z Z_neg VDD VNW pmos_6p0 W=1.22e-06 L=5e-07
.ENDS


.end
