**************************************
* Revision: 1.0
**************************************

*.SCALE METER

.SUBCKT M1_PSUB_CDNS_40254123696109
** N=1781 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_402541236960 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 nmos_5p0 L=6e-07 W=6.81e-06 AD=2.9964e-12 AS=2.9964e-12 PD=1.45e-05 PS=1.45e-05 NRD=0.0646109 NRS=0.0646109 m=1 nf=1 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_402541236962
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_5p0_CDNS_402541236961 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 pmos_5p0 L=6e-07 W=6.81e-06 AD=2.9964e-12 AS=2.9964e-12 PD=1.45e-05 PS=1.45e-05 NRD=0.0646109 NRS=0.0646109 m=1 nf=1 $X=0 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT 018SRAM_cell1_dummy_R
** N=8 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_1 3 4 7 8 9 10
** N=12 EP=6 IP=16 FDC=4
*.SEEDPROM
M0 4 4 7 4 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=3560 $D=8
M1 4 4 9 4 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=4840 $D=8
M2 8 3 4 4 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=3560 $D=8
M3 10 3 4 4 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=4840 $D=8
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 10 12 14 15
** N=19 EP=8 IP=24 FDC=16
*.SEEDPROM
M0 1 3 16 3 nmos_5p0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=180 $Y=7970 $D=2
M1 18 3 1 3 nmos_5p0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=180 $Y=9260 $D=2
M2 3 4 16 3 nmos_5p0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=6340 $D=2
M3 3 4 18 3 nmos_5p0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=10710 $D=2
M4 17 3 3 3 nmos_5p0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=6340 $D=2
M5 19 3 3 3 nmos_5p0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=10710 $D=2
M6 2 3 17 3 nmos_5p0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=2220 $Y=7970 $D=2
M7 19 3 2 3 nmos_5p0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=2220 $Y=9260 $D=2
X8 3 4 10 12 16 17 ICV_1 $T=0 0 0 0 $X=-340 $Y=-340
X9 3 4 18 19 14 15 ICV_1 $T=0 9000 0 0 $X=-340 $Y=8660
.ENDS
***************************************
.SUBCKT 018SRAM_strap1_bndry
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT strapx2b_bndry
** N=10 EP=0 IP=12 FDC=0
.ENDS
***************************************
.SUBCKT dcap_103_novia
** N=2 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT 018SRAM_cell1
** N=8 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT 018SRAM_cell1_2x 1 2 3 5 6 7 8 9 10
** N=12 EP=9 IP=16 FDC=8
*.SEEDPROM
M0 1 5 7 3 nmos_5p0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=180 $Y=3470 $D=2
M1 9 6 1 3 nmos_5p0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=180 $Y=4760 $D=2
M2 3 8 7 3 nmos_5p0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=1840 $D=2
M3 3 10 9 3 nmos_5p0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=6210 $D=2
M4 8 7 3 3 nmos_5p0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=1840 $D=2
M5 10 9 3 3 nmos_5p0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=6210 $D=2
M6 2 5 8 3 nmos_5p0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=2220 $Y=3470 $D=2
M7 10 6 2 3 nmos_5p0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=2220 $Y=4760 $D=2
.ENDS
***************************************
.SUBCKT ICV_3 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
** N=16 EP=15 IP=24 FDC=16
*.SEEDPROM
X0 5 6 2 3 4 9 11 10 12 018SRAM_cell1_2x $T=-3000 0 0 0 $X=-3340 $Y=-340
X1 7 8 2 3 4 13 15 14 16 018SRAM_cell1_2x $T=0 0 0 0 $X=-340 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
** N=26 EP=18 IP=32 FDC=40
*.SEEDPROM
M0 1 20 19 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=8060 $D=8
M1 1 24 23 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=9340 $D=8
M2 20 19 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=8060 $D=8
M3 24 23 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=9340 $D=8
M4 1 22 21 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=8060 $D=8
M5 1 26 25 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=9340 $D=8
M6 22 21 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=8060 $D=8
M7 26 25 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=9340 $D=8
X8 2 3 4 7 8 9 10 11 19 12 20 13 21 14 22 ICV_3 $T=0 0 0 0 $X=-3340 $Y=-340
X9 2 5 6 7 8 9 10 23 15 24 16 25 17 26 18 ICV_3 $T=0 9000 0 0 $X=-3340 $Y=8660
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
** N=30 EP=30 IP=36 FDC=80
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 15 16 17 18 19 20 21 22 ICV_4 $T=-6000 0 0 0 $X=-9340 $Y=-340
X1 1 2 3 4 5 6 11 12 13 14 23 24 25 26 27 28 29 30 ICV_4 $T=0 0 0 0 $X=-3340 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34
** N=50 EP=34 IP=60 FDC=176
*.SEEDPROM
M0 1 36 35 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-8370 $Y=17060 $D=8
M1 1 44 43 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-8370 $Y=18340 $D=8
M2 36 35 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-7230 $Y=17060 $D=8
M3 44 43 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-7230 $Y=18340 $D=8
M4 1 38 37 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-5370 $Y=17060 $D=8
M5 1 46 45 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-5370 $Y=18340 $D=8
M6 38 37 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-4230 $Y=17060 $D=8
M7 46 45 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-4230 $Y=18340 $D=8
M8 1 40 39 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=17060 $D=8
M9 1 48 47 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=18340 $D=8
M10 40 39 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=17060 $D=8
M11 48 47 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=18340 $D=8
M12 1 42 41 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=17060 $D=8
M13 1 50 49 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=18340 $D=8
M14 42 41 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=17060 $D=8
M15 50 49 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=18340 $D=8
X16 1 2 3 4 5 6 11 12 13 14 15 16 17 18 19 20 21 22 35 36
+ 37 38 23 24 25 26 39 40 41 42
+ ICV_5 $T=0 0 0 0 $X=-9340 $Y=-340
X17 1 2 7 8 9 10 11 12 13 14 15 16 17 18 43 44 45 46 27 28
+ 29 30 47 48 49 50 31 32 33 34
+ ICV_5 $T=0 18000 0 0 $X=-9340 $Y=17660
.ENDS
***************************************
.SUBCKT 018SRAM_cell1_dummy 1 2 3 4 5 7
** N=9 EP=6 IP=0 FDC=4
*.SEEDPROM
M0 1 7 2 3 nmos_5p0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=180 $Y=260 $D=2
M1 3 5 1 3 nmos_5p0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=1710 $D=2
M2 5 1 3 3 nmos_5p0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=1710 $D=2
M3 5 7 4 3 nmos_5p0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=2220 $Y=260 $D=2
.ENDS
***************************************
.SUBCKT ICV_7 1 3 4 5 6 7 8 9 10 11
** N=15 EP=10 IP=18 FDC=8
*.SEEDPROM
X0 5 4 1 6 7 3 018SRAM_cell1_dummy $T=-3000 0 0 0 $X=-3340 $Y=-340
X1 9 8 1 10 11 3 018SRAM_cell1_dummy $T=0 0 0 0 $X=-340 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_8 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19
** N=27 EP=18 IP=30 FDC=16
*.SEEDPROM
X0 1 3 4 5 6 7 8 9 10 11 ICV_7 $T=-6000 0 0 0 $X=-9340 $Y=-340
X1 1 3 12 13 14 15 16 17 18 19 ICV_7 $T=0 0 0 0 $X=-3340 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_9
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_10
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_11
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT 018SRAM_strap1
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT 018SRAM_strap1_2x
** N=10 EP=0 IP=12 FDC=0
.ENDS
***************************************
.SUBCKT ICV_12
** N=15 EP=0 IP=20 FDC=0
.ENDS
***************************************
.SUBCKT ICV_13 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22
** N=30 EP=18 IP=33 FDC=16
*.SEEDPROM
X0 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 ICV_8 $T=-3000 0 0 0 $X=-12340 $Y=-340
.ENDS
***************************************
.SUBCKT M1_PSUB$$47122476
** N=5 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pmos_1p2$$46889004 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
X0 1 2 3 4 pmos_5p0_CDNS_402541236961 $T=-155 0 0 0 $X=-1195 $Y=-620
.ENDS
***************************************
.SUBCKT nmos_1p2$$47119404 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
X0 1 2 3 4 nmos_5p0_CDNS_402541236960 $T=-155 0 0 0 $X=-835 $Y=-620
.ENDS
***************************************
.SUBCKT ypass_gate vss 3 b d bb db ypass pcb vdd
** N=26 EP=9 IP=25 FDC=5
*.SEEDPROM
X1 bb b pcb vdd pmos_5p0_CDNS_402541236961 $T=1240 50985 1 0 $X=200 $Y=43555
X2 bb db 3 vdd pmos_5p0_CDNS_402541236961 $T=1250 43050 1 0 $X=210 $Y=35620
X4 b d 3 vdd pmos_1p2$$46889004 $T=1405 15300 1 0 $X=-25 $Y=7790
X5 b d ypass vss nmos_1p2$$47119404 $T=1405 24575 1 0 $X=260 $Y=17090
X6 bb db ypass vss nmos_1p2$$47119404 $T=1405 34595 1 0 $X=260 $Y=27110
.ENDS
***************************************
.SUBCKT mux821 1 2 3 4 5 6 7 8 9 13 14 15 16 17 18 19 20 21 22 23
+ 24 25 26 27 28 29 30 31 32 33 42 43 44 45 46 47 48
** N=86 EP=37 IP=165 FDC=48
*.SEEDPROM
M0 13 42 1 1 nmos_5p0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=1510 $Y=2370 $D=2
M1 16 43 1 1 nmos_5p0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=3750 $Y=2370 $D=2
M2 19 44 1 1 nmos_5p0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=7705 $Y=2370 $D=2
M3 22 45 1 1 nmos_5p0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=9945 $Y=2370 $D=2
M4 25 46 1 1 nmos_5p0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=13895 $Y=2370 $D=2
M5 28 47 1 1 nmos_5p0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=16135 $Y=2370 $D=2
M6 31 48 1 1 nmos_5p0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=20090 $Y=2370 $D=2
M7 2 9 1 1 nmos_5p0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=22330 $Y=2370 $D=2
X9 5 3 7 8 pmos_5p0_CDNS_402541236961 $T=23310 51440 1 0 $X=22270 $Y=44010
X10 5 6 2 8 pmos_5p0_CDNS_402541236961 $T=23320 43505 1 0 $X=22280 $Y=36075
X12 3 4 2 8 pmos_1p2$$46889004 $T=23475 15755 1 0 $X=22045 $Y=8245
X13 3 4 9 1 nmos_1p2$$47119404 $T=23475 25030 1 0 $X=22330 $Y=17545
X14 5 6 9 1 nmos_1p2$$47119404 $T=23475 35050 1 0 $X=22330 $Y=27565
X15 1 13 15 4 14 6 42 7 8 ypass_gate $T=3490 455 1 180 $X=-1160 $Y=0
X16 1 16 18 4 17 6 43 7 8 ypass_gate $T=3490 455 0 0 $X=2385 $Y=0
X17 1 19 21 4 20 6 44 7 8 ypass_gate $T=9685 455 1 180 $X=5035 $Y=0
X18 1 22 24 4 23 6 45 7 8 ypass_gate $T=9685 455 0 0 $X=8580 $Y=0
X19 1 25 27 4 26 6 46 7 8 ypass_gate $T=15875 455 1 180 $X=11225 $Y=0
X20 1 28 30 4 29 6 47 7 8 ypass_gate $T=15875 455 0 0 $X=14770 $Y=0
X21 1 31 33 4 32 6 48 7 8 ypass_gate $T=22070 455 1 180 $X=17420 $Y=0
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_402541236969
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_4025412369640
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_5p0_CDNS_4025412369620
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_4025412369639
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_5p0_CDNS_4025412369629 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pmos_5p0 L=6e-07 W=3.42e-06 AD=8.892e-13 AS=1.5048e-12 PD=4.46e-06 PS=8.6e-06 NRD=0.304094 NRS=0.51462 m=1 nf=2 $X=0 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_402541236968
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_1p2$$202596396
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_5p0_CDNS_4025412369614
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_1p2$$202595372
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$202586156
** N=3 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_5p0_CDNS_4025412369641
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$202587180
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT wen_wm1 vss wep 3 4 5 men 7 8 9 10 11 12 13 14 vdd wen GWEN 18 19
** N=43 EP=19 IP=113 FDC=31
M0 10 wen vss vss nmos_5p0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=1765 $Y=5060 $D=2
M1 7 men vss vss nmos_5p0 L=6e-07 W=1.37e-06 AD=3.562e-13 AS=6.028e-13 PD=1.89e-06 PS=3.62e-06 NRD=0.189781 NRS=0.321168 m=1 nf=1 $X=1765 $Y=8905 $D=2
M2 vss GWEN 10 vss nmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=2885 $Y=5060 $D=2
M3 vss vss 7 vss nmos_5p0 L=6e-07 W=1.37e-06 AD=6.028e-13 AS=3.562e-13 PD=3.62e-06 PS=1.89e-06 NRD=0.321168 NRS=0.189781 m=1 nf=1 $X=2885 $Y=8905 $D=2
M4 3 10 vss vss nmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=5125 $Y=4650 $D=2
M5 11 7 vss vss nmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=5125 $Y=9315 $D=2
M6 4 7 3 vss nmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=7660 $Y=8385 $D=2
M7 8 5 vss vss nmos_5p0 L=6e-07 W=1.37e-06 AD=6.028e-13 AS=6.028e-13 PD=3.62e-06 PS=3.62e-06 NRD=0.321168 NRS=0.321168 m=1 nf=1 $X=8920 $Y=4240 $D=2
M8 12 11 4 vss nmos_5p0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=9970 $Y=9700 $D=2
M9 vss 14 12 vss nmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=11090 $Y=9700 $D=2
M10 vss 4 14 vss nmos_5p0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=13330 $Y=9700 $D=2
M11 13 14 vss vss nmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=14450 $Y=9700 $D=2
M12 wep 8 vss vss nmos_5p0 L=6e-07 W=2.4e-06 AD=7.68e-13 AS=7.68e-13 PD=5.12e-06 PS=5.12e-06 NRD=1.2 NRS=1.2 m=1 nf=3 $X=12720 $Y=4810 $D=2
M13 vss 13 9 vss nmos_5p0 L=6e-07 W=1.37e-06 AD=6.028e-13 AS=6.028e-13 PD=3.62e-06 PS=3.62e-06 NRD=0.321168 NRS=0.321168 m=1 nf=1 $X=17810 $Y=9290 $D=2
M14 men 9 5 vss nmos_5p0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.589e-12 PD=5.58e-06 PS=8.21e-06 NRD=0.229075 NRS=0.30837 m=1 nf=2 $X=20050 $Y=8385 $D=2
M15 vss 13 5 vss nmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=22290 $Y=8385 $D=2
M16 18 wen vdd vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=1765 $Y=600 $D=8
M17 19 men vdd vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=1765 $Y=12055 $D=8
M18 10 GWEN 18 vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=2885 $Y=600 $D=8
M19 7 vss 19 vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=2885 $Y=12055 $D=8
M20 3 10 vdd vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=5125 $Y=600 $D=8
M21 11 7 vdd vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=5125 $Y=12055 $D=8
M22 4 11 3 vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=1.17084e-12 AS=9.988e-13 PD=4.78598e-06 PS=5.42e-06 NRD=0.22722 NRS=0.193833 m=1 nf=1 $X=7660 $Y=12055 $D=8
M23 12 7 4 vdd pmos_5p0 L=6e-07 W=9.6e-07 AD=-6.87097e-13 AS=-6.48697e-13 PD=-2.78573e-06 PS=-2.70573e-06 NRD=-0.745548 NRS=-0.703882 m=1 nf=1 $X=9395 $Y=12055 $D=8
M24 vdd 14 12 vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=1.14386e-12 PD=5.42e-06 PS=4.72975e-06 NRD=0.193833 NRS=0.221983 m=1 nf=1 $X=11090 $Y=12055 $D=8
M25 vdd 4 14 vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=13330 $Y=12055 $D=8
M26 13 14 vdd vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=14450 $Y=12055 $D=8
M27 wep 8 vdd vdd pmos_5p0 L=6e-07 W=6e-06 AD=1.92e-12 AS=1.92e-12 PD=9.92e-06 PS=9.92e-06 NRD=0.48 NRS=0.48 m=1 nf=3 $X=12720 $Y=870 $D=8
M28 men 13 5 vdd pmos_5p0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.58e-06 PS=1.084e-05 NRD=0.229075 NRS=0.387665 m=1 nf=2 $X=20050 $Y=12055 $D=8
X37 vdd 8 5 pmos_5p0_CDNS_4025412369629 $T=8920 2870 1 0 $X=7880 $Y=540
X38 vdd 9 13 pmos_5p0_CDNS_4025412369629 $T=16690 12625 0 0 $X=15650 $Y=12005
.ENDS
***************************************
.SUBCKT M1_PSUB$$44997676
** N=7 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_4025412369612
** N=6 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_4025412369637 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 nmos_5p0 L=6e-07 W=6e-07 AD=2.64e-13 AS=2.64e-13 PD=2.08e-06 PS=2.08e-06 NRD=0.733333 NRS=0.733333 m=1 nf=1 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT pmos_5p0_CDNS_4025412369636
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$46281772
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_4025412369638 1 2 3 4 5
** N=5 EP=5 IP=0 FDC=2
M0 2 4 1 2 nmos_5p0 L=6e-07 W=6e-07 AD=1.56e-13 AS=2.64e-13 PD=1.12e-06 PS=2.08e-06 NRD=0.433333 NRS=0.733333 m=1 nf=1 $X=0 $Y=0 $D=2
M1 3 5 2 2 nmos_5p0 L=6e-07 W=6e-07 AD=2.64e-13 AS=1.56e-13 PD=2.08e-06 PS=1.12e-06 NRD=0.733333 NRS=0.433333 m=1 nf=1 $X=1120 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT pmos_5p0_CDNS_4025412369632 1 2 3 4 5
** N=6 EP=5 IP=0 FDC=2
M0 2 4 1 2 pmos_5p0 L=6e-07 W=1.2e-06 AD=3.12e-13 AS=5.28e-13 PD=1.72e-06 PS=3.28e-06 NRD=0.216667 NRS=0.366667 m=1 nf=1 $X=0 $Y=0 $D=8
M1 3 5 2 2 pmos_5p0 L=6e-07 W=1.2e-06 AD=5.28e-13 AS=3.12e-13 PD=3.28e-06 PS=1.72e-06 NRD=0.366667 NRS=0.216667 m=1 nf=1 $X=1120 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_4025412369633 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 nmos_5p0 L=6e-07 W=1.135e-05 AD=3.3596e-12 AS=3.3596e-12 PD=1.658e-05 PS=1.658e-05 NRD=0.651982 NRS=0.651982 m=1 nf=5 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT pmos_1p2$$46285868
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_5p0_CDNS_4025412369613
** N=6 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$46286892
** N=5 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sacntl_2 vss 2 pcb 4 5 6 7 8 9 10 11 se 19 20 21 22 23 24 25 26
+ 27 vdd men
** N=54 EP=23 IP=83 FDC=39
M0 2 11 vss vss nmos_5p0 L=6e-07 W=2.28e-06 AD=5.928e-13 AS=1.0032e-12 PD=3.32e-06 PS=6.32e-06 NRD=0.45614 NRS=0.77193 m=1 nf=2 $X=795 $Y=26115 $D=2
M1 4 men vss vss nmos_5p0 L=6e-07 W=5.7e-06 AD=1.6872e-12 AS=1.6872e-12 PD=9.8e-06 PS=9.8e-06 NRD=1.29825 NRS=1.29825 m=1 nf=5 $X=855 $Y=4275 $D=2
M2 vss 10 pcb vss nmos_5p0 L=6e-07 W=1.589e-05 AD=4.54e-12 AS=4.54e-12 PD=2.216e-05 PS=2.216e-05 NRD=0.881057 NRS=0.881057 m=1 nf=7 $X=1950 $Y=9235 $D=2
M3 5 4 vss vss nmos_5p0 L=6e-07 W=2.86e-06 AD=7.436e-13 AS=1.2584e-12 PD=3.38e-06 PS=6.6e-06 NRD=0.0909091 NRS=0.153846 m=1 nf=1 $X=10910 $Y=8645 $D=2
M4 6 11 5 vss nmos_5p0 L=6e-07 W=2.86e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=12030 $Y=8645 $D=2
M5 7 27 6 vss nmos_5p0 L=6e-07 W=2.86e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=13150 $Y=8645 $D=2
M6 8 27 7 vss nmos_5p0 L=6e-07 W=2.86e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=14270 $Y=8645 $D=2
M7 9 11 8 vss nmos_5p0 L=6e-07 W=2.86e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=15390 $Y=8645 $D=2
M8 vss 4 9 vss nmos_5p0 L=6e-07 W=2.86e-06 AD=1.2584e-12 AS=7.436e-13 PD=6.6e-06 PS=3.38e-06 NRD=0.153846 NRS=0.0909091 m=1 nf=1 $X=16510 $Y=8645 $D=2
M9 10 7 vss vss nmos_5p0 L=6e-07 W=5.22e-06 AD=1.3572e-12 AS=2.2968e-12 PD=6.26e-06 PS=1.22e-05 NRD=0.199234 NRS=0.337165 m=1 nf=2 $X=18750 $Y=8895 $D=2
M10 11 20 vss vss nmos_5p0 L=6e-07 W=1.44e-06 AD=6.336e-13 AS=6.336e-13 PD=3.76e-06 PS=3.76e-06 NRD=0.305556 NRS=0.305556 m=1 nf=1 $X=21255 $Y=4090 $D=2
M11 se 27 vss vss nmos_5p0 L=6e-07 W=9.08e-06 AD=2.3608e-12 AS=3.178e-12 PD=1.116e-05 PS=1.642e-05 NRD=0.45815 NRS=0.61674 m=1 nf=4 $X=19460 $Y=25030 $D=2
M12 2 11 vdd vdd pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=3.0008e-12 PD=7.86e-06 PS=1.54e-05 NRD=0.152493 NRS=0.258065 m=1 nf=2 $X=795 $Y=20945 $D=8
M13 4 men vdd vdd pmos_5p0 L=6e-07 W=1.135e-05 AD=3.3596e-12 AS=3.3596e-12 PD=1.658e-05 PS=1.658e-05 NRD=0.651982 NRS=0.651982 m=1 nf=5 $X=855 $Y=590 $D=8
M14 27 2 vdd vdd pmos_5p0 L=6e-07 W=6.81e-06 AD=1.7706e-12 AS=2.1792e-12 PD=8.37e-06 PS=1.1e-05 NRD=0.343612 NRS=0.422907 m=1 nf=3 $X=5370 $Y=20990 $D=8
M15 vdd 4 27 vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=8730 $Y=20990 $D=8
M16 pcb 10 vdd vdd pmos_5p0 L=6e-07 W=4.09e-05 AD=1.0634e-11 AS=1.21023e-11 PD=4.61e-05 PS=4.6818e-05 NRD=0.635697 NRS=0.723472 m=1 nf=10 $X=830 $Y=14055 $D=8
M17 7 27 vdd vdd pmos_5p0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.06e-06 PS=9.96e-06 NRD=0.0572687 NRS=0.0969163 m=1 nf=1 $X=14270 $Y=13710 $D=8
M18 vdd 11 7 vdd pmos_5p0 L=6e-07 W=4.54e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=15390 $Y=13710 $D=8
M19 7 4 vdd vdd pmos_5p0 L=6e-07 W=4.54e-06 AD=1.9976e-12 AS=1.1804e-12 PD=9.96e-06 PS=5.06e-06 NRD=0.0969163 NRS=0.0572687 m=1 nf=1 $X=16510 $Y=13710 $D=8
M20 vdd 25 19 vdd pmos_5p0 L=6e-07 W=1.2e-06 AD=5.28e-13 AS=5.28e-13 PD=3.28e-06 PS=3.28e-06 NRD=0.366667 NRS=0.366667 m=1 nf=1 $X=18950 $Y=1670 $D=8
M21 10 7 vdd vdd pmos_5p0 L=6e-07 W=1.362e-05 AD=4.3584e-12 AS=4.3584e-12 PD=2.008e-05 PS=2.008e-05 NRD=0.211454 NRS=0.211454 m=1 nf=3 $X=18750 $Y=13710 $D=8
M22 se 27 vdd vdd pmos_5p0 L=6e-07 W=2.72e-05 AD=7.072e-12 AS=8.0512e-12 PD=3.24e-05 PS=3.856e-05 NRD=0.955882 NRS=1.08824 m=1 nf=10 $X=12740 $Y=20450 $D=8
X23 vdd 11 20 pmos_5p0_CDNS_4025412369629 $T=21255 985 0 0 $X=20215 $Y=365
X27 19 vss 25 vss nmos_5p0_CDNS_4025412369637 $T=18950 4420 0 0 $X=18270 $Y=3800
X31 20 vss 21 4 vss nmos_5p0_CDNS_4025412369638 $T=8080 4420 0 0 $X=7400 $Y=3800
X32 22 vss 23 21 22 nmos_5p0_CDNS_4025412369638 $T=11705 4420 0 0 $X=11025 $Y=3800
X33 24 vss 25 23 24 nmos_5p0_CDNS_4025412369638 $T=15325 4420 0 0 $X=14645 $Y=3800
X34 20 vdd 21 4 vss pmos_5p0_CDNS_4025412369632 $T=8080 1480 0 0 $X=7040 $Y=860
X35 22 vdd 23 21 22 pmos_5p0_CDNS_4025412369632 $T=11705 1480 0 0 $X=10665 $Y=860
X36 24 vdd 25 23 24 pmos_5p0_CDNS_4025412369632 $T=15325 1480 0 0 $X=14285 $Y=860
X37 vss 26 2 vss nmos_5p0_CDNS_4025412369633 $T=5370 25030 0 0 $X=4690 $Y=24410
X38 27 26 4 vss nmos_5p0_CDNS_4025412369633 $T=12415 25030 0 0 $X=11735 $Y=24410
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_4025412369649
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_5p0_CDNS_402541236963
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_5p0_CDNS_4025412369651
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_4025412369644
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT outbuf_oe q vss 3 4 5 15 16 17 18 vdd GWE se qp qn 24
** N=66 EP=15 IP=48 FDC=18
M0 vss 5 q vss nmos_5p0 L=6e-07 W=1.272e-05 AD=3.3072e-12 AS=4.0704e-12 PD=1.584e-05 PS=2.08e-05 NRD=0.735849 NRS=0.90566 m=1 nf=6 $X=395 $Y=2665 $D=2
M1 3 GWE vss vss nmos_5p0 L=6e-07 W=1.6e-06 AD=7.04e-13 AS=7.04e-13 PD=4.08e-06 PS=4.08e-06 NRD=0.275 NRS=0.275 m=1 nf=1 $X=8145 $Y=2720 $D=2
M2 17 3 vss vss nmos_5p0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=9.68e-13 PD=5.28e-06 PS=5.28e-06 NRD=0.2 NRS=0.2 m=1 nf=1 $X=10105 $Y=2700 $D=2
M3 vss 16 4 vss nmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=13175 $Y=12845 $D=2
M4 5 15 4 vss nmos_5p0 L=6e-07 W=6.81e-06 AD=2.1792e-12 AS=2.1792e-12 PD=1.1e-05 PS=1.1e-05 NRD=0.422907 NRS=0.422907 m=1 nf=3 $X=12455 $Y=2720 $D=2
M5 vss se 15 vss nmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=17045 $Y=4035 $D=2
M6 5 qn 18 vss nmos_5p0 L=6e-07 W=5.68e-06 AD=1.4768e-12 AS=1.988e-12 PD=6.72e-06 PS=9.92e-06 NRD=0.183099 NRS=0.246479 m=1 nf=2 $X=19905 $Y=1945 $D=2
M7 vss 3 18 vss nmos_5p0 L=6e-07 W=5.68e-06 AD=1.4768e-12 AS=1.988e-12 PD=6.72e-06 PS=9.92e-06 NRD=0.183099 NRS=0.246479 m=1 nf=2 $X=22145 $Y=1945 $D=2
M8 vdd 5 q vdd pmos_5p0 L=6e-07 W=2.268e-05 AD=5.8968e-12 AS=7.2576e-12 PD=2.58e-05 PS=3.408e-05 NRD=0.412698 NRS=0.507937 m=1 nf=6 $X=395 $Y=6190 $D=8
M9 3 GWE vdd vdd pmos_5p0 L=6e-07 W=4e-06 AD=1.76e-12 AS=1.76e-12 PD=8.88e-06 PS=8.88e-06 NRD=0.11 NRS=0.11 m=1 nf=1 $X=8145 $Y=6395 $D=8
M10 17 3 vdd vdd pmos_5p0 L=6e-07 W=4.5e-06 AD=1.98e-12 AS=1.98e-12 PD=9.88e-06 PS=9.88e-06 NRD=0.0977778 NRS=0.0977778 m=1 nf=1 $X=10105 $Y=6175 $D=8
M11 4 16 vdd vdd pmos_5p0 L=6e-07 W=2.28e-06 AD=5.928e-13 AS=1.24202e-12 PD=3.32e-06 PS=5.60564e-06 NRD=0.45614 NRS=0.955691 m=1 nf=2 $X=12055 $Y=10310 $D=8
M12 5 se 4 vdd pmos_5p0 L=6e-07 W=6.81e-06 AD=2.1792e-12 AS=2.1792e-12 PD=1.1e-05 PS=1.1e-05 NRD=0.422907 NRS=0.422907 m=1 nf=3 $X=12455 $Y=6395 $D=8
M13 16 5 vdd vdd pmos_5p0 L=6e-07 W=1.2e-06 AD=5.28e-13 AS=7.79385e-13 PD=3.28e-06 PS=2.57436e-06 NRD=0.366667 NRS=0.541239 m=1 nf=1 $X=15085 $Y=10250 $D=8
M14 vdd se 15 vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=17045 $Y=7030 $D=8
M15 5 qp 24 vdd pmos_5p0 L=6e-07 W=1.134e-05 AD=2.9484e-12 AS=3.969e-12 PD=1.238e-05 PS=1.841e-05 NRD=0.0917108 NRS=0.123457 m=1 nf=2 $X=19680 $Y=6685 $D=8
M16 vdd 17 24 vdd pmos_5p0 L=6e-07 W=1.134e-05 AD=2.9484e-12 AS=3.969e-12 PD=1.238e-05 PS=1.841e-05 NRD=0.0917108 NRS=0.123457 m=1 nf=2 $X=21920 $Y=6685 $D=8
X20 vss 16 5 vss nmos_5p0_CDNS_4025412369637 $T=15150 13365 1 0 $X=14470 $Y=12145
.ENDS
***************************************
.SUBCKT M1_NWELL_CDNS_4025412369636
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_4025412369611 1 2 3 4 5 6
** N=6 EP=6 IP=0 FDC=2
M0 2 4 1 6 nmos_5p0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=0 $Y=0 $D=2
M1 3 5 2 6 nmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=1120 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT nmos_1p2$$46883884 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 nmos_5p0 L=6e-07 W=1.134e-05 AD=4.9896e-12 AS=4.9896e-12 PD=2.356e-05 PS=2.356e-05 NRD=0.0388007 NRS=0.0388007 m=1 nf=1 $X=-155 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT nmos_1p2$$46563372 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
M0 2 3 1 4 nmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=-155 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT pmos_5p0_CDNS_402541236966 1 2 3 4 5 6
** N=6 EP=6 IP=0 FDC=2
M0 2 4 1 6 pmos_5p0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=0 $Y=0 $D=8
M1 3 5 2 6 pmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=1120 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT pmos_1p2$$46273580 1 2 3
** N=3 EP=3 IP=3 FDC=1
M0 2 3 1 1 pmos_5p0 L=6e-07 W=2.28e-06 AD=5.928e-13 AS=1.0032e-12 PD=3.32e-06 PS=6.32e-06 NRD=0.45614 NRS=0.77193 m=1 nf=2 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT pmos_1p2$$46887980 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pmos_5p0 L=6e-07 W=1.361e-05 AD=5.9884e-12 AS=5.9884e-12 PD=2.81e-05 PS=2.81e-05 NRD=0.0323292 NRS=0.0323292 m=1 nf=1 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT din vss 2 3 4 5 6 7 8 d db 11 12 vdd datain men wep
** N=69 EP=16 IP=73 FDC=24
M0 2 4 vss vss nmos_5p0 L=6e-07 W=1.361e-05 AD=5.9884e-12 AS=5.9884e-12 PD=2.81e-05 PS=2.81e-05 NRD=0.0323292 NRS=0.0323292 m=1 nf=1 $X=260 $Y=10430 $D=2
M1 3 wep vss vss nmos_5p0 L=6e-07 W=1.14e-06 AD=7.866e-13 AS=7.923e-13 PD=3.66e-06 PS=3.67e-06 NRD=0.605263 NRS=0.609649 m=1 nf=1 $X=3600 $Y=38320 $D=2
M2 vss 7 4 vss nmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=11165 $Y=8655 $D=2
M3 3 wep vdd vdd pmos_5p0 L=6e-07 W=2.97e-06 AD=1.13602e-12 AS=1.7523e-12 PD=4.5e-06 PS=8.3e-06 NRD=0.515152 NRS=0.794613 m=1 nf=2 $X=3025 $Y=35440 $D=8
M4 vdd 2 11 vdd pmos_5p0 L=6e-07 W=1.134e-05 AD=4.9896e-12 AS=4.9896e-12 PD=2.356e-05 PS=2.356e-05 NRD=0.0388007 NRS=0.0388007 m=1 nf=1 $X=6980 $Y=26220 $D=8
X5 4 vdd 7 vdd pmos_5p0_CDNS_402541236961 $T=11165 455 0 0 $X=10125 $Y=-165
X6 d 2 3 vdd pmos_1p2$$46889004 $T=2655 26220 0 0 $X=1225 $Y=25510
X7 db 11 3 vdd pmos_1p2$$46889004 $T=4895 26220 0 0 $X=3465 $Y=25510
X10 5 vss 6 datain 5 vss nmos_5p0_CDNS_4025412369611 $T=2765 1790 1 0 $X=2085 $Y=210
X11 6 7 8 12 men vss nmos_5p0_CDNS_4025412369611 $T=6905 725 0 0 $X=6225 $Y=105
X12 d 2 wep vss nmos_1p2$$46883884 $T=2655 12695 0 0 $X=1510 $Y=12010
X13 db 11 wep vss nmos_1p2$$46883884 $T=4895 12695 0 0 $X=3750 $Y=12010
X14 11 vss 2 vss nmos_1p2$$46883884 $T=7135 12695 0 0 $X=5990 $Y=12010
X15 vss 12 men vss nmos_1p2$$46563372 $T=3470 9035 0 0 $X=2325 $Y=8350
X16 vss 8 4 vss nmos_1p2$$46563372 $T=7060 10495 1 0 $X=5915 $Y=8860
X17 5 vdd 6 datain 5 vdd pmos_5p0_CDNS_402541236966 $T=2765 3195 0 0 $X=1725 $Y=2575
X18 6 7 8 men 12 vdd pmos_5p0_CDNS_402541236966 $T=6905 3605 0 0 $X=5865 $Y=2985
X19 vdd 12 men pmos_1p2$$46273580 $T=2920 7175 1 0 $X=1490 $Y=5355
X20 vdd 8 4 pmos_1p2$$46273580 $T=7060 8140 1 0 $X=5630 $Y=6320
X21 vdd 2 4 pmos_1p2$$46887980 $T=415 26220 0 0 $X=-1015 $Y=25510
.ENDS
***************************************
.SUBCKT nmos_1p2$$46553132
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$46897196 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
M0 2 3 1 4 pmos_5p0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.58e-06 PS=1.084e-05 NRD=0.229075 NRS=0.387665 m=1 nf=2 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT pmos_1p2$$46898220
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_1p2$$46551084
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sa 1 vss 3 4 qn qp 7 pcb vdd d db se
** N=105 EP=12 IP=47 FDC=27
M0 1 vss vss vss nmos_5p0 L=6e-07 W=3.41e-06 AD=8.866e-13 AS=1.5004e-12 PD=3.93e-06 PS=7.7e-06 NRD=0.0762463 NRS=0.129032 m=1 nf=1 $X=11660 $Y=16585 $D=2
M1 3 4 1 vss nmos_5p0 L=6e-07 W=3.41e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=12780 $Y=16585 $D=2
M2 4 1 3 vss nmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=1.7732e-12 PD=7.86e-06 PS=7.86e-06 NRD=0.152493 NRS=0.152493 m=1 nf=2 $X=13900 $Y=16585 $D=2
M3 7 4 vss vss nmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=15170 $Y=8510 $D=2
M4 1 4 3 vss nmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=1.7732e-12 PD=7.86e-06 PS=7.86e-06 NRD=0.152493 NRS=0.152493 m=1 nf=2 $X=16140 $Y=16585 $D=2
M5 4 1 3 vss nmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=1.7732e-12 PD=7.86e-06 PS=7.86e-06 NRD=0.152493 NRS=0.152493 m=1 nf=2 $X=18380 $Y=16585 $D=2
M6 vss 7 qp vss nmos_5p0 L=6e-07 W=6.81e-06 AD=1.7706e-12 AS=2.1792e-12 PD=8.37e-06 PS=1.1e-05 NRD=0.343612 NRS=0.422907 m=1 nf=3 $X=17410 $Y=8510 $D=2
M7 1 4 3 vss nmos_5p0 L=6e-07 W=3.41e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=20620 $Y=16585 $D=2
M8 qn 1 vss vss nmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=20770 $Y=8510 $D=2
M9 3 se vss vss nmos_5p0 L=6e-07 W=2.272e-05 AD=5.9072e-12 AS=6.9296e-12 PD=2.688e-05 PS=3.328e-05 NRD=0.732394 NRS=0.859155 m=1 nf=8 $X=12945 $Y=12550 $D=2
M10 vss vss 1 vss nmos_5p0 L=6e-07 W=3.41e-06 AD=1.5004e-12 AS=8.866e-13 PD=7.7e-06 PS=3.93e-06 NRD=0.129032 NRS=0.0762463 m=1 nf=1 $X=21740 $Y=16585 $D=2
M11 4 vdd vdd vdd pmos_5p0 L=6e-07 W=9.1e-07 AD=2.366e-13 AS=4.004e-13 PD=1.43e-06 PS=2.7e-06 NRD=0.285714 NRS=0.483516 m=1 nf=1 $X=13985 $Y=24010 $D=8
M12 vdd 1 4 vdd pmos_5p0 L=6e-07 W=9.1e-07 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=15105 $Y=24010 $D=8
M13 d pcb vdd vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=15755 $Y=30660 $D=8
M14 7 4 vdd vdd pmos_5p0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.589e-12 PD=5.58e-06 PS=8.21e-06 NRD=0.229075 NRS=0.30837 m=1 nf=2 $X=15170 $Y=4385 $D=8
M15 4 pcb 1 vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=16875 $Y=26330 $D=8
M16 db pcb d vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=16875 $Y=30660 $D=8
M17 1 4 vdd vdd pmos_5p0 L=6e-07 W=1.82e-06 AD=4.732e-13 AS=4.732e-13 PD=2.86e-06 PS=2.86e-06 NRD=0.571429 NRS=0.571429 m=1 nf=2 $X=16225 $Y=24010 $D=8
M18 vdd pcb db vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=17995 $Y=30660 $D=8
M19 4 1 vdd vdd pmos_5p0 L=6e-07 W=9.1e-07 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=18465 $Y=24010 $D=8
M20 qp 7 vdd vdd pmos_5p0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.1804e-12 PD=5.58e-06 PS=5.58e-06 NRD=0.229075 NRS=0.229075 m=1 nf=2 $X=17410 $Y=4385 $D=8
M21 vdd vdd 4 vdd pmos_5p0 L=6e-07 W=9.1e-07 AD=4.004e-13 AS=2.366e-13 PD=2.7e-06 PS=1.43e-06 NRD=0.483516 NRS=0.285714 m=1 nf=1 $X=19585 $Y=24010 $D=8
M22 qn 1 vdd vdd pmos_5p0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.589e-12 PD=5.58e-06 PS=8.21e-06 NRD=0.229075 NRS=0.30837 m=1 nf=2 $X=19650 $Y=4385 $D=8
X28 db 1 se vdd pmos_1p2$$46897196 $T=12475 26330 0 0 $X=11045 $Y=25620
X29 d 4 se vdd pmos_1p2$$46897196 $T=12475 30660 0 0 $X=11045 $Y=29950
X30 d 4 se vdd pmos_1p2$$46897196 $T=20400 26330 0 0 $X=18970 $Y=25620
X31 db 1 se vdd pmos_1p2$$46897196 $T=20400 30660 0 0 $X=18970 $Y=29950
.ENDS
***************************************
.SUBCKT saout_R_m2 1 vss q pcb datain men vdd b[7] bb[7] WEN b[0] bb[0] bb[1] b[1] b[2] bb[2] bb[3] b[3] b[4] bb[4]
+ bb[5] b[5] b[6] bb[6] 54 ypass[0] ypass[1] ypass[2] GWE ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] GWEN 74 75 76 77 78
+ 79 80
** N=131 EP=42 IP=161 FDC=187
*.SEEDPROM
X0 vss 54 b[7] 70 bb[7] 73 pcb vdd ypass[7] 74 bb[0] b[0] 75 bb[1] b[1] 76 bb[2] b[2] 77 bb[3]
+ b[3] 78 bb[4] b[4] 79 bb[5] b[5] 80 bb[6] b[6] ypass[0] ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6]
+ mux821 $T=2765 83310 0 0 $X=-1345 $Y=83305
X1 vss 1 85 87 93 men 83 88 92 82 86 89 91 90 vdd WEN GWEN 81 84 wen_wm1 $T=1610 -16880 0 0 $X=100 $Y=-17420
X2 vss 94 pcb 68 99 100 101 102 104 107 108 72 106 97 71 98 69 103 105 96
+ 95 vdd men
+ sacntl_2 $T=3160 115 0 0 $X=425 $Y=-5
X3 q vss 109 111 112 114 113 110 116 vdd GWE 72 130 131 115 outbuf_oe $T=3160 27545 0 0 $X=500 $Y=25750
X4 vss 117 120 125 118 121 123 124 70 73 122 119 vdd datain men 1 din $T=1615 39025 0 0 $X=500 $Y=38740
X5 126 vss 128 127 131 130 129 pcb vdd 70 73 72 sa $T=3160 43040 0 0 $X=1375 $Y=42060
.ENDS
***************************************
.SUBCKT ICV_14 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
** N=16 EP=15 IP=24 FDC=16
*.SEEDPROM
X0 5 6 2 3 4 9 11 10 12 018SRAM_cell1_2x $T=0 0 0 0 $X=-340 $Y=-340
X1 7 8 2 3 4 13 15 14 16 018SRAM_cell1_2x $T=3000 0 0 0 $X=2660 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_15 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
** N=26 EP=18 IP=32 FDC=40
*.SEEDPROM
M0 1 20 19 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=8060 $D=8
M1 1 24 23 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=9340 $D=8
M2 20 19 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=8060 $D=8
M3 24 23 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=9340 $D=8
M4 1 22 21 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=8060 $D=8
M5 1 26 25 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=9340 $D=8
M6 22 21 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=8060 $D=8
M7 26 25 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=9340 $D=8
X8 2 3 4 7 8 9 10 11 19 12 20 13 21 14 22 ICV_14 $T=0 0 0 0 $X=-340 $Y=-340
X9 2 5 6 7 8 9 10 23 15 24 16 25 17 26 18 ICV_14 $T=0 9000 0 0 $X=-340 $Y=8660
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
** N=30 EP=30 IP=36 FDC=80
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 15 16 17 18 19 20 21 22 ICV_15 $T=0 0 0 0 $X=-340 $Y=-340
X1 1 2 3 4 5 6 11 12 13 14 23 24 25 26 27 28 29 30 ICV_15 $T=6000 0 0 0 $X=5660 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_17 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34
** N=50 EP=34 IP=60 FDC=176
*.SEEDPROM
M0 1 36 35 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=17060 $D=8
M1 1 44 43 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=18340 $D=8
M2 36 35 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=17060 $D=8
M3 44 43 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=18340 $D=8
M4 1 38 37 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=17060 $D=8
M5 1 46 45 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=18340 $D=8
M6 38 37 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=17060 $D=8
M7 46 45 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=18340 $D=8
M8 1 40 39 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=6630 $Y=17060 $D=8
M9 1 48 47 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=6630 $Y=18340 $D=8
M10 40 39 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=7770 $Y=17060 $D=8
M11 48 47 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=7770 $Y=18340 $D=8
M12 1 42 41 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=9630 $Y=17060 $D=8
M13 1 50 49 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=9630 $Y=18340 $D=8
M14 42 41 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=10770 $Y=17060 $D=8
M15 50 49 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=10770 $Y=18340 $D=8
X16 1 2 3 4 5 6 11 12 13 14 15 16 17 18 19 20 21 22 35 36
+ 37 38 23 24 25 26 39 40 41 42
+ ICV_16 $T=0 0 0 0 $X=-340 $Y=-340
X17 1 2 7 8 9 10 11 12 13 14 15 16 17 18 43 44 45 46 27 28
+ 29 30 47 48 49 50 31 32 33 34
+ ICV_16 $T=0 18000 0 0 $X=-340 $Y=17660
.ENDS
***************************************
.SUBCKT new_dummyrow_unit 7 9 43 45 47 49 51 53 55 57 59 61 63 65 67 69 71 73 75 77
+ 79 81 83 85 87 89 91 93 95 97 99 101 103 105
** N=105 EP=34 IP=120 FDC=64
*.SEEDPROM
X0 7 9 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 ICV_8 $T=3310 885 1 180 $X=-30 $Y=545
X1 7 9 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 ICV_8 $T=15310 885 1 180 $X=11970 $Y=545
X2 7 9 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 ICV_8 $T=30310 885 1 180 $X=26970 $Y=545
X3 7 9 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 ICV_8 $T=42310 885 1 180 $X=38970 $Y=545
.ENDS
***************************************
.SUBCKT saout_m2 1 VSS q datain pcb men VDD b[0] bb[0] WEN b[7] bb[7] bb[6] b[6] b[5] bb[5] bb[4] b[4] b[3] bb[3]
+ bb[2] b[2] b[1] bb[1] 54 ypass[7] ypass[6] ypass[5] GWE ypass[4] ypass[3] ypass[2] ypass[1] ypass[0] GWEN 78 79 80 81 82
+ 83 84
** N=135 EP=42 IP=161 FDC=187
*.SEEDPROM
X0 VSS 54 b[0] 74 bb[0] 77 pcb VDD ypass[0] 78 bb[7] b[7] 79 bb[6] b[6] 80 bb[5] b[5] 81 bb[4]
+ b[4] 82 bb[3] b[3] 83 bb[2] b[2] 84 bb[1] b[1] ypass[7] ypass[6] ypass[5] ypass[4] ypass[3] ypass[2] ypass[1]
+ mux821 $T=2765 83345 0 0 $X=-1345 $Y=83340
X1 VSS 1 89 91 97 men 87 92 96 86 90 93 95 94 VDD WEN GWEN 85 88 wen_wm1 $T=1610 -16845 0 0 $X=100 $Y=-17385
X2 VSS 98 pcb 72 103 104 105 106 108 111 112 76 110 101 75 102 73 107 109 100
+ 99 VDD men
+ sacntl_2 $T=3160 150 0 0 $X=425 $Y=30
X3 q VSS 113 115 116 118 117 114 120 VDD GWE 76 134 135 119 outbuf_oe $T=3160 27580 0 0 $X=500 $Y=25785
X4 VSS 121 124 129 122 125 127 128 74 77 126 123 VDD datain men 1 din $T=1615 39060 0 0 $X=500 $Y=38775
X5 130 VSS 132 131 135 134 133 pcb VDD 74 77 76 sa $T=3160 43075 0 0 $X=1375 $Y=42095
.ENDS
***************************************
.SUBCKT ICV_18 8 11 12 13 14 15 16
** N=16 EP=7 IP=22 FDC=8
*.SEEDPROM
X1 11 12 8 8 8 13 15 14 16 018SRAM_cell1_2x $T=0 0 0 0 $X=-340 $Y=-340
.ENDS
***************************************
.SUBCKT rcol4_64 VSS tblhl pcb[4] VDD DWL WEN[6] pcb[6] 8 9 men WEN[4] 12 13 WEN[7] pcb[7] 16 17 WEN[5] pcb[5] 20
+ 21 WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] GWE GWEN ypass[1] ypass[0] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] din[5]
+ q[5] din[7] q[7] din[4] q[4] din[6] q[6] 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445
** N=665 EP=103 IP=1279 FDC=2834
*.SEEDPROM
M0 195 VSS 83 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=1715 $Y=151295 $D=2
M1 83 VSS 197 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=1715 $Y=195005 $D=2
M2 VSS 194 195 VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=2165 $Y=152745 $D=2
M3 VSS 196 197 VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=2165 $Y=193375 $D=2
M4 194 195 VSS VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=3305 $Y=152745 $D=2
M5 196 197 VSS VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=3305 $Y=193375 $D=2
M6 194 VSS 82 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=3755 $Y=151295 $D=2
M7 82 VSS 196 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=3755 $Y=195005 $D=2
M8 450 VSS 61 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=115715 $Y=151295 $D=2
M9 61 VSS 452 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=115715 $Y=168005 $D=2
M10 454 VSS 61 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=115715 $Y=169295 $D=2
M11 61 DWL 456 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=115715 $Y=186005 $D=2
M12 446 DWL 61 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=115715 $Y=187295 $D=2
M13 61 DWL 448 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=115715 $Y=195005 $D=2
M14 VSS VDD 450 VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=116165 $Y=152745 $D=2
M15 VSS VDD 452 VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=116165 $Y=166375 $D=2
M16 VSS VDD 454 VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=116165 $Y=170745 $D=2
M17 VSS VDD 456 VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=116165 $Y=184375 $D=2
M18 VSS VDD 446 VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=116165 $Y=188745 $D=2
M19 VSS VDD 448 VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=116165 $Y=193375 $D=2
M20 451 VSS VSS VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=117305 $Y=152745 $D=2
M21 453 VSS VSS VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=117305 $Y=166375 $D=2
M22 455 VSS VSS VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=117305 $Y=170745 $D=2
M23 457 VSS VSS VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=117305 $Y=184375 $D=2
M24 447 VSS VSS VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=117305 $Y=188745 $D=2
M25 449 VSS VSS VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=117305 $Y=193375 $D=2
M26 55 61 VSS VSS nmos_5p0 L=6e-07 W=2.76e-06 AD=7.176e-13 AS=1.2144e-12 PD=3.8e-06 PS=7.28e-06 NRD=0.376812 NRS=0.637681 m=1 nf=2 $X=116215 $Y=69445 $D=2
M27 tblhl 55 VSS VSS nmos_5p0 L=6e-07 W=1.7e-05 AD=4.42e-12 AS=7.48e-12 PD=1.804e-05 PS=3.576e-05 NRD=0.0611765 NRS=0.103529 m=1 nf=2 $X=116235 $Y=54020 $D=2
M28 63 VDD VSS VSS nmos_5p0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=5.016e-13 PD=2.18e-06 PS=4.04e-06 NRD=0.912281 NRS=1.54386 m=1 nf=2 $X=116460 $Y=85710 $D=2
M29 451 VSS 62 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=117755 $Y=151295 $D=2
M30 62 VSS 453 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=117755 $Y=168005 $D=2
M31 455 VSS 62 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=117755 $Y=169295 $D=2
M32 62 DWL 457 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=117755 $Y=186005 $D=2
M33 447 DWL 62 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=117755 $Y=187295 $D=2
M34 62 DWL 449 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=117755 $Y=195005 $D=2
M35 VDD 194 195 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=2165 $Y=154595 $D=8
M36 VDD 650 652 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=2165 $Y=155875 $D=8
M37 VDD 651 653 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=2165 $Y=163595 $D=8
M38 VDD 654 656 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=2165 $Y=164875 $D=8
M39 VDD 655 657 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=2165 $Y=172595 $D=8
M40 VDD 658 660 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=2165 $Y=173875 $D=8
M41 VDD 659 661 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=2165 $Y=181595 $D=8
M42 VDD 662 664 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=2165 $Y=182875 $D=8
M43 VDD 663 665 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=2165 $Y=190595 $D=8
M44 VDD 196 197 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=2165 $Y=191875 $D=8
M45 194 195 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=3305 $Y=154595 $D=8
M46 650 652 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=3305 $Y=155875 $D=8
M47 651 653 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=3305 $Y=163595 $D=8
M48 654 656 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=3305 $Y=164875 $D=8
M49 655 657 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=3305 $Y=172595 $D=8
M50 658 660 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=3305 $Y=173875 $D=8
M51 659 661 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=3305 $Y=181595 $D=8
M52 662 664 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=3305 $Y=182875 $D=8
M53 663 665 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=3305 $Y=190595 $D=8
M54 196 197 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=3305 $Y=191875 $D=8
M55 VDD 323 325 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=8165 $Y=154595 $D=8
M56 VDD 541 540 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=8165 $Y=155875 $D=8
M57 VDD 549 548 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=8165 $Y=190595 $D=8
M58 VDD 243 245 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=8165 $Y=191875 $D=8
M59 323 325 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=9305 $Y=154595 $D=8
M60 541 540 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=9305 $Y=155875 $D=8
M61 549 548 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=9305 $Y=190595 $D=8
M62 243 245 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=9305 $Y=191875 $D=8
M63 636 ypass[7] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=9160 $Y=87735 $D=8
M64 VDD 319 321 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=11165 $Y=154595 $D=8
M65 VDD 543 542 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=11165 $Y=155875 $D=8
M66 VDD 551 550 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=11165 $Y=190595 $D=8
M67 VDD 239 241 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=11165 $Y=191875 $D=8
M68 319 321 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=12305 $Y=154595 $D=8
M69 543 542 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=12305 $Y=155875 $D=8
M70 551 550 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=12305 $Y=190595 $D=8
M71 239 241 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=12305 $Y=191875 $D=8
M72 637 ypass[6] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=11690 $Y=87735 $D=8
M73 VDD 315 317 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=14165 $Y=154595 $D=8
M74 VDD 545 544 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=14165 $Y=155875 $D=8
M75 VDD 553 552 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=14165 $Y=190595 $D=8
M76 VDD 235 237 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=14165 $Y=191875 $D=8
M77 315 317 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=15305 $Y=154595 $D=8
M78 545 544 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=15305 $Y=155875 $D=8
M79 553 552 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=15305 $Y=190595 $D=8
M80 235 237 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=15305 $Y=191875 $D=8
M81 638 ypass[5] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=15355 $Y=87735 $D=8
M82 VDD 311 313 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=17165 $Y=154595 $D=8
M83 VDD 547 546 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=17165 $Y=155875 $D=8
M84 VDD 555 554 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=17165 $Y=190595 $D=8
M85 VDD 231 233 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=17165 $Y=191875 $D=8
M86 311 313 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=18305 $Y=154595 $D=8
M87 547 546 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=18305 $Y=155875 $D=8
M88 555 554 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=18305 $Y=190595 $D=8
M89 231 233 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=18305 $Y=191875 $D=8
M90 639 ypass[4] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=17885 $Y=87735 $D=8
M91 VDD 203 205 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=20165 $Y=154595 $D=8
M92 VDD 557 556 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=20165 $Y=155875 $D=8
M93 VDD 565 564 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=20165 $Y=190595 $D=8
M94 VDD 259 261 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=20165 $Y=191875 $D=8
M95 203 205 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=21305 $Y=154595 $D=8
M96 557 556 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=21305 $Y=155875 $D=8
M97 565 564 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=21305 $Y=190595 $D=8
M98 259 261 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=21305 $Y=191875 $D=8
M99 640 ypass[3] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=21545 $Y=87735 $D=8
M100 VDD 199 201 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=23165 $Y=154595 $D=8
M101 VDD 559 558 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=23165 $Y=155875 $D=8
M102 VDD 567 566 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=23165 $Y=190595 $D=8
M103 VDD 255 257 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=23165 $Y=191875 $D=8
M104 199 201 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=24305 $Y=154595 $D=8
M105 559 558 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=24305 $Y=155875 $D=8
M106 567 566 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=24305 $Y=190595 $D=8
M107 255 257 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=24305 $Y=191875 $D=8
M108 641 ypass[2] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=24075 $Y=87735 $D=8
M109 VDD 211 213 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=26165 $Y=154595 $D=8
M110 VDD 561 560 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=26165 $Y=155875 $D=8
M111 VDD 569 568 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=26165 $Y=190595 $D=8
M112 VDD 251 253 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=26165 $Y=191875 $D=8
M113 211 213 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=27305 $Y=154595 $D=8
M114 561 560 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=27305 $Y=155875 $D=8
M115 569 568 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=27305 $Y=190595 $D=8
M116 251 253 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=27305 $Y=191875 $D=8
M117 642 ypass[1] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=27740 $Y=87735 $D=8
M118 VDD 207 209 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=29165 $Y=154595 $D=8
M119 VDD 563 562 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=29165 $Y=155875 $D=8
M120 VDD 571 570 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=29165 $Y=190595 $D=8
M121 VDD 247 249 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=29165 $Y=191875 $D=8
M122 207 209 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=30305 $Y=154595 $D=8
M123 563 562 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=30305 $Y=155875 $D=8
M124 571 570 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=30305 $Y=190595 $D=8
M125 247 249 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=30305 $Y=191875 $D=8
M126 460 ypass[0] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=30270 $Y=87735 $D=8
M127 VDD 339 341 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=35165 $Y=154595 $D=8
M128 VDD 468 469 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=35165 $Y=155875 $D=8
M129 VDD 476 477 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=35165 $Y=190595 $D=8
M130 VDD 355 357 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=35165 $Y=191875 $D=8
M131 458 ypass[7] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=33945 $Y=87735 $D=8
M132 339 341 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=36305 $Y=154595 $D=8
M133 468 469 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=36305 $Y=155875 $D=8
M134 476 477 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=36305 $Y=190595 $D=8
M135 355 357 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=36305 $Y=191875 $D=8
M136 532 ypass[6] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=36470 $Y=87735 $D=8
M137 VDD 335 337 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=38165 $Y=154595 $D=8
M138 VDD 466 467 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=38165 $Y=155875 $D=8
M139 VDD 474 475 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=38165 $Y=190595 $D=8
M140 VDD 351 353 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=38165 $Y=191875 $D=8
M141 335 337 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=39305 $Y=154595 $D=8
M142 466 467 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=39305 $Y=155875 $D=8
M143 474 475 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=39305 $Y=190595 $D=8
M144 351 353 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=39305 $Y=191875 $D=8
M145 VDD 331 333 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=41165 $Y=154595 $D=8
M146 VDD 464 465 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=41165 $Y=155875 $D=8
M147 VDD 472 473 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=41165 $Y=190595 $D=8
M148 VDD 347 349 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=41165 $Y=191875 $D=8
M149 531 ypass[5] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=40135 $Y=87735 $D=8
M150 331 333 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=42305 $Y=154595 $D=8
M151 464 465 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=42305 $Y=155875 $D=8
M152 472 473 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=42305 $Y=190595 $D=8
M153 347 349 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=42305 $Y=191875 $D=8
M154 530 ypass[4] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=42665 $Y=87735 $D=8
M155 VDD 327 329 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=44165 $Y=154595 $D=8
M156 VDD 462 463 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=44165 $Y=155875 $D=8
M157 VDD 470 471 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=44165 $Y=190595 $D=8
M158 VDD 343 345 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=44165 $Y=191875 $D=8
M159 327 329 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=45305 $Y=154595 $D=8
M160 462 463 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=45305 $Y=155875 $D=8
M161 470 471 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=45305 $Y=190595 $D=8
M162 343 345 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=45305 $Y=191875 $D=8
M163 VDD 275 277 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=47165 $Y=154595 $D=8
M164 VDD 484 485 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=47165 $Y=155875 $D=8
M165 VDD 492 493 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=47165 $Y=190595 $D=8
M166 VDD 291 293 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=47165 $Y=191875 $D=8
M167 529 ypass[3] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=46325 $Y=87735 $D=8
M168 275 277 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=48305 $Y=154595 $D=8
M169 484 485 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=48305 $Y=155875 $D=8
M170 492 493 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=48305 $Y=190595 $D=8
M171 291 293 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=48305 $Y=191875 $D=8
M172 528 ypass[2] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=48855 $Y=87735 $D=8
M173 VDD 271 273 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=50165 $Y=154595 $D=8
M174 VDD 482 483 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=50165 $Y=155875 $D=8
M175 VDD 490 491 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=50165 $Y=190595 $D=8
M176 VDD 287 289 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=50165 $Y=191875 $D=8
M177 271 273 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=51305 $Y=154595 $D=8
M178 482 483 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=51305 $Y=155875 $D=8
M179 490 491 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=51305 $Y=190595 $D=8
M180 287 289 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=51305 $Y=191875 $D=8
M181 VDD 267 269 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=53165 $Y=154595 $D=8
M182 VDD 480 481 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=53165 $Y=155875 $D=8
M183 VDD 488 489 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=53165 $Y=190595 $D=8
M184 VDD 283 285 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=53165 $Y=191875 $D=8
M185 527 ypass[1] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=52520 $Y=87735 $D=8
M186 267 269 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=54305 $Y=154595 $D=8
M187 480 481 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=54305 $Y=155875 $D=8
M188 488 489 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=54305 $Y=190595 $D=8
M189 283 285 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=54305 $Y=191875 $D=8
M190 VDD 263 265 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=56165 $Y=154595 $D=8
M191 VDD 478 479 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=56165 $Y=155875 $D=8
M192 VDD 486 487 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=56165 $Y=190595 $D=8
M193 VDD 279 281 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=56165 $Y=191875 $D=8
M194 526 ypass[0] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=55050 $Y=87735 $D=8
M195 263 265 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=57305 $Y=154595 $D=8
M196 478 479 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=57305 $Y=155875 $D=8
M197 486 487 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=57305 $Y=190595 $D=8
M198 279 281 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=57305 $Y=191875 $D=8
M199 VDD 371 373 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=62165 $Y=154595 $D=8
M200 VDD 573 572 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=62165 $Y=155875 $D=8
M201 VDD 581 580 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=62165 $Y=190595 $D=8
M202 VDD 610 611 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=62165 $Y=191875 $D=8
M203 371 373 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=63305 $Y=154595 $D=8
M204 573 572 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=63305 $Y=155875 $D=8
M205 581 580 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=63305 $Y=190595 $D=8
M206 610 611 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=63305 $Y=191875 $D=8
M207 643 ypass[7] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=63160 $Y=87735 $D=8
M208 VDD 367 369 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=65165 $Y=154595 $D=8
M209 VDD 575 574 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=65165 $Y=155875 $D=8
M210 VDD 583 582 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=65165 $Y=190595 $D=8
M211 VDD 608 609 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=65165 $Y=191875 $D=8
M212 367 369 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=66305 $Y=154595 $D=8
M213 575 574 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=66305 $Y=155875 $D=8
M214 583 582 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=66305 $Y=190595 $D=8
M215 608 609 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=66305 $Y=191875 $D=8
M216 644 ypass[6] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=65690 $Y=87735 $D=8
M217 VDD 363 365 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=68165 $Y=154595 $D=8
M218 VDD 577 576 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=68165 $Y=155875 $D=8
M219 VDD 585 584 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=68165 $Y=190595 $D=8
M220 VDD 606 607 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=68165 $Y=191875 $D=8
M221 363 365 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=69305 $Y=154595 $D=8
M222 577 576 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=69305 $Y=155875 $D=8
M223 585 584 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=69305 $Y=190595 $D=8
M224 606 607 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=69305 $Y=191875 $D=8
M225 645 ypass[5] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=69355 $Y=87735 $D=8
M226 VDD 359 361 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=71165 $Y=154595 $D=8
M227 VDD 579 578 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=71165 $Y=155875 $D=8
M228 VDD 587 586 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=71165 $Y=190595 $D=8
M229 VDD 604 605 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=71165 $Y=191875 $D=8
M230 359 361 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=72305 $Y=154595 $D=8
M231 579 578 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=72305 $Y=155875 $D=8
M232 587 586 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=72305 $Y=190595 $D=8
M233 604 605 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=72305 $Y=191875 $D=8
M234 646 ypass[4] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=71885 $Y=87735 $D=8
M235 VDD 219 221 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=74165 $Y=154595 $D=8
M236 VDD 589 588 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=74165 $Y=155875 $D=8
M237 VDD 597 596 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=74165 $Y=190595 $D=8
M238 VDD 618 619 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=74165 $Y=191875 $D=8
M239 219 221 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=75305 $Y=154595 $D=8
M240 589 588 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=75305 $Y=155875 $D=8
M241 597 596 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=75305 $Y=190595 $D=8
M242 618 619 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=75305 $Y=191875 $D=8
M243 647 ypass[3] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=75545 $Y=87735 $D=8
M244 VDD 215 217 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=77165 $Y=154595 $D=8
M245 VDD 591 590 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=77165 $Y=155875 $D=8
M246 VDD 599 598 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=77165 $Y=190595 $D=8
M247 VDD 616 617 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=77165 $Y=191875 $D=8
M248 215 217 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=78305 $Y=154595 $D=8
M249 591 590 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=78305 $Y=155875 $D=8
M250 599 598 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=78305 $Y=190595 $D=8
M251 616 617 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=78305 $Y=191875 $D=8
M252 648 ypass[2] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=78075 $Y=87735 $D=8
M253 VDD 227 229 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=80165 $Y=154595 $D=8
M254 VDD 593 592 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=80165 $Y=155875 $D=8
M255 VDD 601 600 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=80165 $Y=190595 $D=8
M256 VDD 614 615 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=80165 $Y=191875 $D=8
M257 227 229 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=81305 $Y=154595 $D=8
M258 593 592 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=81305 $Y=155875 $D=8
M259 601 600 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=81305 $Y=190595 $D=8
M260 614 615 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=81305 $Y=191875 $D=8
M261 649 ypass[1] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=81740 $Y=87735 $D=8
M262 VDD 223 225 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=83165 $Y=154595 $D=8
M263 VDD 595 594 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=83165 $Y=155875 $D=8
M264 VDD 603 602 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=83165 $Y=190595 $D=8
M265 VDD 612 613 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=83165 $Y=191875 $D=8
M266 223 225 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=84305 $Y=154595 $D=8
M267 595 594 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=84305 $Y=155875 $D=8
M268 603 602 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=84305 $Y=190595 $D=8
M269 612 613 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=84305 $Y=191875 $D=8
M270 461 ypass[0] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=84270 $Y=87735 $D=8
M271 VDD 387 389 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=89165 $Y=154595 $D=8
M272 VDD 500 501 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=89165 $Y=155875 $D=8
M273 VDD 508 509 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=89165 $Y=190595 $D=8
M274 VDD 626 627 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=89165 $Y=191875 $D=8
M275 459 ypass[7] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=87945 $Y=87735 $D=8
M276 387 389 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=90305 $Y=154595 $D=8
M277 500 501 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=90305 $Y=155875 $D=8
M278 508 509 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=90305 $Y=190595 $D=8
M279 626 627 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=90305 $Y=191875 $D=8
M280 539 ypass[6] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=90470 $Y=87735 $D=8
M281 VDD 383 385 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=92165 $Y=154595 $D=8
M282 VDD 498 499 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=92165 $Y=155875 $D=8
M283 VDD 506 507 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=92165 $Y=190595 $D=8
M284 VDD 624 625 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=92165 $Y=191875 $D=8
M285 383 385 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=93305 $Y=154595 $D=8
M286 498 499 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=93305 $Y=155875 $D=8
M287 506 507 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=93305 $Y=190595 $D=8
M288 624 625 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=93305 $Y=191875 $D=8
M289 VDD 379 381 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=95165 $Y=154595 $D=8
M290 VDD 496 497 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=95165 $Y=155875 $D=8
M291 VDD 504 505 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=95165 $Y=190595 $D=8
M292 VDD 622 623 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=95165 $Y=191875 $D=8
M293 538 ypass[5] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=94135 $Y=87735 $D=8
M294 379 381 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=96305 $Y=154595 $D=8
M295 496 497 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=96305 $Y=155875 $D=8
M296 504 505 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=96305 $Y=190595 $D=8
M297 622 623 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=96305 $Y=191875 $D=8
M298 537 ypass[4] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=96665 $Y=87735 $D=8
M299 VDD 375 377 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=98165 $Y=154595 $D=8
M300 VDD 494 495 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=98165 $Y=155875 $D=8
M301 VDD 502 503 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=98165 $Y=190595 $D=8
M302 VDD 620 621 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=98165 $Y=191875 $D=8
M303 375 377 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=99305 $Y=154595 $D=8
M304 494 495 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=99305 $Y=155875 $D=8
M305 502 503 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=99305 $Y=190595 $D=8
M306 620 621 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=99305 $Y=191875 $D=8
M307 VDD 307 309 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=101165 $Y=154595 $D=8
M308 VDD 516 517 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=101165 $Y=155875 $D=8
M309 VDD 524 525 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=101165 $Y=190595 $D=8
M310 VDD 634 635 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=101165 $Y=191875 $D=8
M311 536 ypass[3] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=100325 $Y=87735 $D=8
M312 307 309 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=102305 $Y=154595 $D=8
M313 516 517 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=102305 $Y=155875 $D=8
M314 524 525 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=102305 $Y=190595 $D=8
M315 634 635 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=102305 $Y=191875 $D=8
M316 535 ypass[2] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=102855 $Y=87735 $D=8
M317 VDD 303 305 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=104165 $Y=154595 $D=8
M318 VDD 514 515 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=104165 $Y=155875 $D=8
M319 VDD 522 523 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=104165 $Y=190595 $D=8
M320 VDD 632 633 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=104165 $Y=191875 $D=8
M321 303 305 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=105305 $Y=154595 $D=8
M322 514 515 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=105305 $Y=155875 $D=8
M323 522 523 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=105305 $Y=190595 $D=8
M324 632 633 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=105305 $Y=191875 $D=8
M325 VDD 299 301 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=107165 $Y=154595 $D=8
M326 VDD 512 513 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=107165 $Y=155875 $D=8
M327 VDD 520 521 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=107165 $Y=190595 $D=8
M328 VDD 630 631 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=107165 $Y=191875 $D=8
M329 534 ypass[1] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=106520 $Y=87735 $D=8
M330 299 301 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=108305 $Y=154595 $D=8
M331 512 513 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=108305 $Y=155875 $D=8
M332 520 521 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=108305 $Y=190595 $D=8
M333 630 631 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=108305 $Y=191875 $D=8
M334 VDD 295 297 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=110165 $Y=154595 $D=8
M335 VDD 510 511 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=110165 $Y=155875 $D=8
M336 VDD 518 519 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=110165 $Y=190595 $D=8
M337 VDD 628 629 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=110165 $Y=191875 $D=8
M338 533 ypass[0] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=109050 $Y=87735 $D=8
M339 295 297 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=111305 $Y=154595 $D=8
M340 510 511 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=111305 $Y=155875 $D=8
M341 518 519 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=111305 $Y=190595 $D=8
M342 628 629 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=111305 $Y=191875 $D=8
M343 VDD VSS VDD VDD pmos_5p0 L=2.365e-06 W=8.19e-05 AD=0 AS=6.1309e-11 PD=0 PS=0.000217698 NRD=0 NRS=11.8457 m=1 nf=36 $X=1805 $Y=145970 $D=8
M344 61 pcb[4] VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=6.35965e-12 PD=7.86e-06 PS=1.737e-05 NRD=0.152493 NRS=0.546921 m=1 nf=2 $X=116100 $Y=135875 $D=8
M345 62 pcb[4] VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=6.35965e-12 PD=7.86e-06 PS=1.737e-05 NRD=0.152493 NRS=0.546921 m=1 nf=2 $X=116100 $Y=139750 $D=8
M346 55 61 VDD VDD pmos_5p0 L=6e-07 W=7.02e-06 AD=1.8252e-12 AS=3.0888e-12 PD=8.06e-06 PS=1.58e-05 NRD=0.148148 NRS=0.250712 m=1 nf=2 $X=116215 $Y=72345 $D=8
M347 tblhl 55 VDD VDD pmos_5p0 L=6e-07 W=2.128e-05 AD=5.5328e-12 AS=9.3632e-12 PD=2.232e-05 PS=4.432e-05 NRD=0.0488722 NRS=0.0827068 m=1 nf=2 $X=116235 $Y=41975 $D=8
M348 63 VDD VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=2.33887e-12 PD=4.29e-06 PS=9.09e-06 NRD=0.444444 NRS=1.06061 m=1 nf=2 $X=116315 $Y=87735 $D=8
X349 61 61 VDD VSS nmos_5p0_CDNS_402541236960 $T=117260 108370 0 180 $X=115980 $Y=100940
X350 62 62 VDD VSS nmos_5p0_CDNS_402541236960 $T=117260 118390 0 180 $X=115980 $Y=110960
X352 61 61 63 VDD pmos_5p0_CDNS_402541236961 $T=117260 99095 0 180 $X=115620 $Y=91665
X353 62 62 63 VDD pmos_5p0_CDNS_402541236961 $T=117260 126845 0 180 $X=115620 $Y=119415
X354 62 61 pcb[4] VDD pmos_5p0_CDNS_402541236961 $T=117270 134780 0 180 $X=115630 $Y=127350
X355 VSS VDD 446 447 448 449 ICV_1 $T=115535 187035 0 0 $X=115195 $Y=186695
X356 61 62 VSS VDD 450 451 452 453 ICV_2 $T=115535 151035 0 0 $X=115195 $Y=150695
X357 61 62 VSS VDD 454 455 456 457 ICV_2 $T=115535 169035 0 0 $X=115195 $Y=168695
X368 VDD VSS WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] 390 391 392 393 394 395 9 8 462 463
+ 464 465 466 467 468 469 470 471 472 473 474 475 476 477
+ ICV_6 $T=37535 155535 1 180 $X=34195 $Y=155195
X369 VDD VSS WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] 396 397 398 399 400 401 402 403 478 479
+ 480 481 482 483 484 485 486 487 488 489 490 491 492 493
+ ICV_6 $T=49535 155535 1 180 $X=46195 $Y=155195
X370 VDD VSS WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] 404 405 406 407 408 409 13 12 494 495
+ 496 497 498 499 500 501 502 503 504 505 506 507 508 509
+ ICV_6 $T=91535 155535 1 180 $X=88195 $Y=155195
X371 VDD VSS WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] 410 411 412 413 414 415 416 417 510 511
+ 512 513 514 515 516 517 518 519 520 521 522 523 524 525
+ ICV_6 $T=103535 155535 1 180 $X=100195 $Y=155195
X372 VSS VSS 198 199 200 201 202 203 204 205 ICV_7 $T=22535 151035 1 180 $X=19195 $Y=150695
X373 VSS VSS 206 207 208 209 210 211 212 213 ICV_7 $T=28535 151035 1 180 $X=25195 $Y=150695
X374 VSS VSS 214 215 216 217 218 219 220 221 ICV_7 $T=76535 151035 1 180 $X=73195 $Y=150695
X375 VSS VSS 222 223 224 225 226 227 228 229 ICV_7 $T=82535 151035 1 180 $X=79195 $Y=150695
X376 VSS DWL 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 ICV_8 $T=10535 196035 0 180 $X=7195 $Y=191195
X377 VSS DWL 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261 ICV_8 $T=22535 196035 0 180 $X=19195 $Y=191195
X378 VSS VSS 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 ICV_8 $T=49535 151035 1 180 $X=46195 $Y=150695
X379 VSS DWL 278 279 280 281 282 283 284 285 286 287 288 289 290 291 292 293 ICV_8 $T=49535 196035 0 180 $X=46195 $Y=191195
X380 VSS VSS 294 295 296 297 298 299 300 301 302 303 304 305 306 307 308 309 ICV_8 $T=103535 151035 1 180 $X=100195 $Y=150695
X395 VSS VSS 310 311 312 313 314 315 316 317 318 319 320 321 322 323 324 325 ICV_13 $T=7535 151035 1 180 $X=4195 $Y=150695
X396 VSS VSS 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 ICV_13 $T=34535 151035 1 180 $X=31195 $Y=150695
X397 VSS DWL 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 ICV_13 $T=34535 196035 0 180 $X=31195 $Y=191195
X398 VSS VSS 358 359 360 361 362 363 364 365 366 367 368 369 370 371 372 373 ICV_13 $T=61535 151035 1 180 $X=58195 $Y=150695
X399 VSS VSS 374 375 376 377 378 379 380 381 382 383 384 385 386 387 388 389 ICV_13 $T=88535 151035 1 180 $X=85195 $Y=150695
X400 153 VSS q[5] pcb[6] din[5] men VDD 8 9 WEN[6] 396 397 398 399 400 401 402 403 390 391
+ 392 393 394 395 458 ypass[0] ypass[1] ypass[2] GWE ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] GWEN 526 527 528 529 530
+ 531 532
+ saout_R_m2 $T=60970 30 1 180 $X=22805 $Y=-18280
X401 154 VSS q[7] pcb[4] din[7] men VDD 12 13 WEN[4] 410 411 412 413 414 415 416 417 404 405
+ 406 407 408 409 459 ypass[0] ypass[1] ypass[2] GWE ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] GWEN 533 534 535 536 537
+ 538 539
+ saout_R_m2 $T=114970 30 1 180 $X=76805 $Y=-18280
X402 VDD VSS WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] 437 436 435 434 433 432 431 430 540 541
+ 542 543 544 545 546 547 548 549 550 551 552 553 554 555
+ ICV_17 $T=7535 155535 0 0 $X=7195 $Y=155195
X403 VDD VSS WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] 421 420 419 418 423 422 17 16 556 557
+ 558 559 560 561 562 563 564 565 566 567 568 569 570 571
+ ICV_17 $T=19535 155535 0 0 $X=19195 $Y=155195
X404 VDD VSS WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] 445 444 443 442 441 440 439 438 572 573
+ 574 575 576 577 578 579 580 581 582 583 584 585 586 587
+ ICV_17 $T=61535 155535 0 0 $X=61195 $Y=155195
X405 VDD VSS WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] 427 426 425 424 429 428 21 20 588 589
+ 590 591 592 593 594 595 596 597 598 599 600 601 602 603
+ ICV_17 $T=73535 155535 0 0 $X=73195 $Y=155195
X406 VSS DWL 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621
+ 622 623 624 625 626 627 628 629 630 631 632 633 634 635
+ new_dummyrow_unit $T=61225 196920 1 0 $X=61195 $Y=191195
X407 155 VSS q[4] din[4] pcb[7] men VDD 16 17 WEN[7] 437 436 435 434 433 432 431 430 421 420
+ 419 418 423 422 460 ypass[7] ypass[6] ypass[5] GWE ypass[4] ypass[3] ypass[2] ypass[1] ypass[0] GWEN 636 637 638 639 640
+ 641 642
+ saout_m2 $T=5100 -5 0 0 $X=3755 $Y=-17780
X408 156 VSS q[6] din[6] pcb[5] men VDD 20 21 WEN[5] 445 444 443 442 441 440 439 438 427 426
+ 425 424 429 428 461 ypass[7] ypass[6] ypass[5] GWE ypass[4] ypass[3] ypass[2] ypass[1] ypass[0] GWEN 643 644 645 646 647
+ 648 649
+ saout_m2 $T=59100 -5 0 0 $X=57755 $Y=-17780
X409 VSS 82 83 650 651 652 653 ICV_18 $T=4535 155535 1 180 $X=1195 $Y=155195
X410 VSS 82 83 654 655 656 657 ICV_18 $T=4535 164535 1 180 $X=1195 $Y=164195
X411 VSS 82 83 658 659 660 661 ICV_18 $T=4535 173535 1 180 $X=1195 $Y=173195
X412 VSS 82 83 662 663 664 665 ICV_18 $T=4535 182535 1 180 $X=1195 $Y=182195
.ENDS
***************************************
.SUBCKT M1_PSUB_CDNS_402541236962
** N=666 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pmos_1p2$$47815724
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_19
** N=4 EP=0 IP=8 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$48624684
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT M1_PSUB_CDNS_4025412369620
** N=1201 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_4025412369694 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nmos_5p0 L=1.2e-06 W=6e-07 AD=2.64e-13 AS=2.64e-13 PD=2.08e-06 PS=2.08e-06 NRD=0.733333 NRS=0.733333 m=1 nf=1 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT pmos_5p0_CDNS_4025412369691 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pmos_5p0 L=1.2e-06 W=9e-07 AD=3.96e-13 AS=3.96e-13 PD=2.68e-06 PS=2.68e-06 NRD=0.488889 NRS=0.488889 m=1 nf=1 $X=0 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nmos_1p2$$47342636
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$47512620
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$47513644
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_4025412369660
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_1p2$$47514668
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT xpredec1_xa
** N=29 EP=0 IP=36 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$47330348_161 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
M0 2 3 1 4 pmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT alatch vss ab a vdd enb en
** N=16 EP=6 IP=24 FDC=8
M0 ab 11 vss vss nmos_5p0 L=6e-07 W=3.64e-06 AD=9.464e-13 AS=1.6016e-12 PD=4.68e-06 PS=9.04e-06 NRD=0.285714 NRS=0.483516 m=1 nf=2 $X=2590 $Y=1475 $D=2
M1 vss ab 12 vss nmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=3710 $Y=12935 $D=2
M2 a en 11 vss nmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=6280 $Y=1020 $D=2
M3 12 enb 11 vss nmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=6280 $Y=12935 $D=2
M4 ab 11 vdd vdd pmos_5p0 L=6e-07 W=9.08e-06 AD=2.3608e-12 AS=3.9952e-12 PD=1.012e-05 PS=1.992e-05 NRD=0.114537 NRS=0.193833 m=1 nf=2 $X=2590 $Y=4695 $D=8
M5 a enb 11 vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=6280 $Y=5895 $D=8
X10 12 vdd ab vdd pmos_1p2$$47330348_161 $T=3865 11540 1 0 $X=2435 $Y=9910
X11 11 12 en vdd pmos_1p2$$47330348_161 $T=6435 11540 1 0 $X=5005 $Y=9910
.ENDS
***************************************
.SUBCKT M1_PSUB$$47335468
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pmos_1p2$$47337516 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pmos_5p0 L=6e-07 W=1.633e-05 AD=7.1852e-12 AS=7.1852e-12 PD=3.354e-05 PS=3.354e-05 NRD=0.0269443 NRS=0.0269443 m=1 nf=1 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nmos_1p2$$47336492 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nmos_5p0 L=6e-07 W=6.58e-06 AD=2.8952e-12 AS=2.8952e-12 PD=1.404e-05 PS=1.404e-05 NRD=0.0668693 NRS=0.0668693 m=1 nf=1 $X=-155 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT xpredec1_bot 1 2 3 10 11 12 13
** N=32 EP=7 IP=19 FDC=12
X0 1 32 11 10 13 12 alatch $T=350 -3160 0 0 $X=-100 $Y=-3165
X2 10 2 32 pmos_1p2$$47337516 $T=3910 18340 0 0 $X=2480 $Y=17635
X3 10 3 2 pmos_1p2$$47337516 $T=6480 18340 0 0 $X=5050 $Y=17635
X4 1 2 32 nmos_1p2$$47336492 $T=3910 36070 0 0 $X=2765 $Y=35385
X5 1 3 2 nmos_1p2$$47336492 $T=6480 36070 0 0 $X=5335 $Y=35385
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_4025412369666
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$47109164 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 pmos_5p0 L=6e-07 W=3.42e-06 AD=8.892e-13 AS=1.5048e-12 PD=4.46e-06 PS=8.6e-06 NRD=0.304094 NRS=0.51462 m=1 nf=2 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT xpredec1 vss men vdd clk A[2] A[1] A[0] x[7] x[6] x[5] x[4] x[3] x[2] x[1] x[0]
** N=91 EP=15 IP=199 FDC=108
M0 77 18 51 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=3.2435e-12 AS=7.36025e-12 PD=1.2995e-05 PS=2.613e-05 NRD=0.0208417 NRS=0.0472946 m=1 nf=1 $X=1700 $Y=2310 $D=2
M1 76 19 77 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=2820 $Y=2310 $D=2
M2 vss 20 76 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=3940 $Y=2310 $D=2
M3 vss 51 x[7] vss nmos_5p0 L=6e-07 W=1.362e-05 AD=3.5412e-12 AS=4.3584e-12 PD=1.518e-05 PS=2.008e-05 NRD=0.171806 NRS=0.211454 m=1 nf=3 $X=1700 $Y=48000 $D=2
M4 78 21 vss vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=5060 $Y=2310 $D=2
M5 79 19 78 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=6180 $Y=2310 $D=2
M6 54 18 79 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=7.36025e-12 AS=3.2435e-12 PD=2.613e-05 PS=1.2995e-05 NRD=0.0472946 NRS=0.0208417 m=1 nf=1 $X=7300 $Y=2310 $D=2
M7 x[6] 54 vss vss nmos_5p0 L=6e-07 W=1.362e-05 AD=4.3584e-12 AS=3.5412e-12 PD=2.008e-05 PS=1.518e-05 NRD=0.211454 NRS=0.171806 m=1 nf=3 $X=5060 $Y=48000 $D=2
M8 81 18 57 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=3.2435e-12 AS=7.36025e-12 PD=1.2995e-05 PS=2.613e-05 NRD=0.0208417 NRS=0.0472946 m=1 nf=1 $X=9870 $Y=2310 $D=2
M9 80 22 81 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=10990 $Y=2310 $D=2
M10 vss 20 80 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=12110 $Y=2310 $D=2
M11 vss 57 x[5] vss nmos_5p0 L=6e-07 W=1.362e-05 AD=3.5412e-12 AS=4.3584e-12 PD=1.518e-05 PS=2.008e-05 NRD=0.171806 NRS=0.211454 m=1 nf=3 $X=9870 $Y=48000 $D=2
M12 82 21 vss vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=13230 $Y=2310 $D=2
M13 83 22 82 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=14350 $Y=2310 $D=2
M14 60 18 83 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=7.36025e-12 AS=3.2435e-12 PD=2.613e-05 PS=1.2995e-05 NRD=0.0472946 NRS=0.0208417 m=1 nf=1 $X=15470 $Y=2310 $D=2
M15 x[4] 60 vss vss nmos_5p0 L=6e-07 W=1.362e-05 AD=4.3584e-12 AS=3.5412e-12 PD=2.008e-05 PS=1.518e-05 NRD=0.211454 NRS=0.171806 m=1 nf=3 $X=13230 $Y=48000 $D=2
M16 85 23 63 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=3.2435e-12 AS=7.36025e-12 PD=1.2995e-05 PS=2.613e-05 NRD=0.0208417 NRS=0.0472946 m=1 nf=1 $X=18035 $Y=2310 $D=2
M17 84 19 85 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=19155 $Y=2310 $D=2
M18 vss 20 84 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=20275 $Y=2310 $D=2
M19 vss 63 x[3] vss nmos_5p0 L=6e-07 W=1.362e-05 AD=3.5412e-12 AS=4.3584e-12 PD=1.518e-05 PS=2.008e-05 NRD=0.171806 NRS=0.211454 m=1 nf=3 $X=18035 $Y=48000 $D=2
M20 86 21 vss vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=21395 $Y=2310 $D=2
M21 87 19 86 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=22515 $Y=2310 $D=2
M22 66 23 87 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=7.36025e-12 AS=3.2435e-12 PD=2.613e-05 PS=1.2995e-05 NRD=0.0472946 NRS=0.0208417 m=1 nf=1 $X=23635 $Y=2310 $D=2
M23 x[2] 66 vss vss nmos_5p0 L=6e-07 W=1.362e-05 AD=4.3584e-12 AS=3.5412e-12 PD=2.008e-05 PS=1.518e-05 NRD=0.211454 NRS=0.171806 m=1 nf=3 $X=21395 $Y=48000 $D=2
M24 89 23 69 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=3.2435e-12 AS=7.36025e-12 PD=1.2995e-05 PS=2.613e-05 NRD=0.0208417 NRS=0.0472946 m=1 nf=1 $X=26205 $Y=2310 $D=2
M25 88 22 89 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=27325 $Y=2310 $D=2
M26 vss 20 88 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=28445 $Y=2310 $D=2
M27 vss 69 x[1] vss nmos_5p0 L=6e-07 W=1.362e-05 AD=3.5412e-12 AS=4.3584e-12 PD=1.518e-05 PS=2.008e-05 NRD=0.171806 NRS=0.211454 m=1 nf=3 $X=26205 $Y=48000 $D=2
M28 90 21 vss vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=29565 $Y=2310 $D=2
M29 91 22 90 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=30685 $Y=2310 $D=2
M30 72 23 91 vss nmos_5p0 L=6e-07 W=1.2475e-05 AD=7.36025e-12 AS=3.2435e-12 PD=2.613e-05 PS=1.2995e-05 NRD=0.0472946 NRS=0.0208417 m=1 nf=1 $X=31805 $Y=2310 $D=2
M31 x[0] 72 vss vss nmos_5p0 L=6e-07 W=1.362e-05 AD=4.3584e-12 AS=3.5412e-12 PD=2.008e-05 PS=1.518e-05 NRD=0.211454 NRS=0.171806 m=1 nf=3 $X=29565 $Y=48000 $D=2
M32 17 men vss vss nmos_5p0 L=6e-07 W=1.91e-06 AD=4.966e-13 AS=8.404e-13 PD=2.43e-06 PS=4.7e-06 NRD=0.136126 NRS=0.230366 m=1 nf=1 $X=37165 $Y=51200 $D=2
M33 vss clk 17 vss nmos_5p0 L=6e-07 W=1.91e-06 AD=8.404e-13 AS=4.966e-13 PD=4.7e-06 PS=2.43e-06 NRD=0.230366 NRS=0.136126 m=1 nf=1 $X=38285 $Y=51200 $D=2
M34 vss 17 16 vss nmos_5p0 L=6e-07 W=1.36e-06 AD=5.984e-13 AS=5.984e-13 PD=3.6e-06 PS=3.6e-06 NRD=0.323529 NRS=0.323529 m=1 nf=1 $X=45140 $Y=51180 $D=2
M35 vdd 18 51 vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=2.7118e-12 AS=4.5892e-12 PD=1.095e-05 PS=2.174e-05 NRD=0.0249281 NRS=0.042186 m=1 nf=1 $X=1700 $Y=21650 $D=8
M36 51 19 vdd vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=2820 $Y=21650 $D=8
M37 vdd 20 51 vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=3940 $Y=21650 $D=8
M38 vdd 51 x[7] vdd pmos_5p0 L=6e-07 W=3.402e-05 AD=8.8452e-12 AS=1.08864e-11 PD=3.558e-05 PS=4.728e-05 NRD=0.0687831 NRS=0.0846561 m=1 nf=3 $X=1700 $Y=35260 $D=8
M39 54 21 vdd vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=5060 $Y=21650 $D=8
M40 vdd 19 54 vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=6180 $Y=21650 $D=8
M41 54 18 vdd vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=4.5892e-12 AS=2.7118e-12 PD=2.174e-05 PS=1.095e-05 NRD=0.042186 NRS=0.0249281 m=1 nf=1 $X=7300 $Y=21650 $D=8
M42 x[6] 54 vdd vdd pmos_5p0 L=6e-07 W=3.402e-05 AD=1.08864e-11 AS=8.8452e-12 PD=4.728e-05 PS=3.558e-05 NRD=0.0846561 NRS=0.0687831 m=1 nf=3 $X=5060 $Y=35260 $D=8
M43 vdd 18 57 vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=2.7118e-12 AS=4.5892e-12 PD=1.095e-05 PS=2.174e-05 NRD=0.0249281 NRS=0.042186 m=1 nf=1 $X=9870 $Y=21650 $D=8
M44 57 22 vdd vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=10990 $Y=21650 $D=8
M45 vdd 20 57 vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=12110 $Y=21650 $D=8
M46 vdd 57 x[5] vdd pmos_5p0 L=6e-07 W=3.402e-05 AD=8.8452e-12 AS=1.08864e-11 PD=3.558e-05 PS=4.728e-05 NRD=0.0687831 NRS=0.0846561 m=1 nf=3 $X=9870 $Y=35260 $D=8
M47 60 21 vdd vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=13230 $Y=21650 $D=8
M48 vdd 22 60 vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=14350 $Y=21650 $D=8
M49 60 18 vdd vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=4.5892e-12 AS=2.7118e-12 PD=2.174e-05 PS=1.095e-05 NRD=0.042186 NRS=0.0249281 m=1 nf=1 $X=15470 $Y=21650 $D=8
M50 x[4] 60 vdd vdd pmos_5p0 L=6e-07 W=3.402e-05 AD=1.08864e-11 AS=8.8452e-12 PD=4.728e-05 PS=3.558e-05 NRD=0.0846561 NRS=0.0687831 m=1 nf=3 $X=13230 $Y=35260 $D=8
M51 vdd 23 63 vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=2.7118e-12 AS=4.5892e-12 PD=1.095e-05 PS=2.174e-05 NRD=0.0249281 NRS=0.042186 m=1 nf=1 $X=18035 $Y=21650 $D=8
M52 63 19 vdd vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=19155 $Y=21650 $D=8
M53 vdd 20 63 vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=20275 $Y=21650 $D=8
M54 vdd 63 x[3] vdd pmos_5p0 L=6e-07 W=3.402e-05 AD=8.8452e-12 AS=1.08864e-11 PD=3.558e-05 PS=4.728e-05 NRD=0.0687831 NRS=0.0846561 m=1 nf=3 $X=18035 $Y=35260 $D=8
M55 66 21 vdd vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=21395 $Y=21650 $D=8
M56 vdd 19 66 vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=22515 $Y=21650 $D=8
M57 66 23 vdd vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=4.5892e-12 AS=2.7118e-12 PD=2.174e-05 PS=1.095e-05 NRD=0.042186 NRS=0.0249281 m=1 nf=1 $X=23635 $Y=21650 $D=8
M58 x[2] 66 vdd vdd pmos_5p0 L=6e-07 W=3.402e-05 AD=1.08864e-11 AS=8.8452e-12 PD=4.728e-05 PS=3.558e-05 NRD=0.0846561 NRS=0.0687831 m=1 nf=3 $X=21395 $Y=35260 $D=8
M59 vdd 23 69 vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=2.7118e-12 AS=4.5892e-12 PD=1.095e-05 PS=2.174e-05 NRD=0.0249281 NRS=0.042186 m=1 nf=1 $X=26205 $Y=21650 $D=8
M60 69 22 vdd vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=27325 $Y=21650 $D=8
M61 vdd 20 69 vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=28445 $Y=21650 $D=8
M62 vdd 69 x[1] vdd pmos_5p0 L=6e-07 W=3.402e-05 AD=8.8452e-12 AS=1.08864e-11 PD=3.558e-05 PS=4.728e-05 NRD=0.0687831 NRS=0.0846561 m=1 nf=3 $X=26205 $Y=35260 $D=8
M63 72 21 vdd vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=29565 $Y=21650 $D=8
M64 vdd 22 72 vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=30685 $Y=21650 $D=8
M65 72 23 vdd vdd pmos_5p0 L=6e-07 W=1.043e-05 AD=4.5892e-12 AS=2.7118e-12 PD=2.174e-05 PS=1.095e-05 NRD=0.042186 NRS=0.0249281 m=1 nf=1 $X=31805 $Y=21650 $D=8
M66 x[0] 72 vdd vdd pmos_5p0 L=6e-07 W=3.402e-05 AD=1.08864e-11 AS=8.8452e-12 PD=4.728e-05 PS=3.558e-05 NRD=0.0846561 NRS=0.0687831 m=1 nf=3 $X=29565 $Y=35260 $D=8
M67 74 men vdd vdd pmos_5p0 L=6e-07 W=2.275e-06 AD=5.915e-13 AS=1.35362e-12 PD=2.795e-06 PS=5.74e-06 NRD=0.114286 NRS=0.261538 m=1 nf=1 $X=37165 $Y=47525 $D=8
M68 17 clk 74 vdd pmos_5p0 L=6e-07 W=2.275e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=38285 $Y=47525 $D=8
M69 75 clk 17 vdd pmos_5p0 L=6e-07 W=2.275e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=39405 $Y=47525 $D=8
M70 vdd men 75 vdd pmos_5p0 L=6e-07 W=2.275e-06 AD=1.35362e-12 AS=5.915e-13 PD=5.74e-06 PS=2.795e-06 NRD=0.261538 NRS=0.114286 m=1 nf=1 $X=40525 $Y=47525 $D=8
X80 vss 18 23 vdd A[2] 17 16 xpredec1_bot $T=34205 3160 0 0 $X=33675 $Y=-5
X81 vss 19 22 vdd A[1] 17 16 xpredec1_bot $T=42655 3160 0 0 $X=42125 $Y=-5
X82 vss 20 21 vdd A[0] 17 16 xpredec1_bot $T=51110 3160 0 0 $X=50580 $Y=-5
X85 vdd 16 17 pmos_1p2$$47109164 $T=44700 47595 0 0 $X=42105 $Y=46910
.ENDS
***************************************
.SUBCKT M1_PACTIVE_CDNS_4025412369671
** N=7 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_4025412369678 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nmos_5p0 L=6e-07 W=1.92e-05 AD=4.992e-12 AS=5.6832e-12 PD=2.44e-05 PS=2.896e-05 NRD=1.35417 NRS=1.54167 m=1 nf=10 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT pmos_5p0_CDNS_4025412369680 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pmos_5p0 L=6e-07 W=4.72e-05 AD=1.2272e-11 AS=1.39712e-11 PD=5.24e-05 PS=6.256e-05 NRD=0.550847 NRS=0.627119 m=1 nf=10 $X=0 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT wen_v2 vss 2 vdd wen clk IGWEN GWE
** N=50 EP=7 IP=93 FDC=30
M0 vss wen 29 vss nmos_5p0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=2545 $Y=1065 $D=2
M1 12 wen vss vss nmos_5p0 L=6e-07 W=6e-06 AD=1.92e-12 AS=1.92e-12 PD=9.92e-06 PS=9.92e-06 NRD=0.48 NRS=0.48 m=1 nf=3 $X=1260 $Y=16070 $D=2
M2 32 clk vss vss nmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=3665 $Y=1065 $D=2
M3 2 32 vss vss nmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=5905 $Y=1475 $D=2
M4 30 32 29 vss nmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=8440 $Y=545 $D=2
M5 34 2 30 vss nmos_5p0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=10750 $Y=1860 $D=2
M6 vss 35 34 vss nmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=11870 $Y=1860 $D=2
M7 vss 30 35 vss nmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=14110 $Y=1860 $D=2
M8 16 35 vss vss nmos_5p0 L=6e-07 W=2.4e-06 AD=6.24e-13 AS=1.056e-12 PD=3.44e-06 PS=6.56e-06 NRD=0.433333 NRS=0.733333 m=1 nf=2 $X=16465 $Y=1620 $D=2
M9 16 2 31 vss nmos_5p0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.58e-06 PS=1.084e-05 NRD=0.229075 NRS=0.387665 m=1 nf=2 $X=19750 $Y=545 $D=2
M10 33 32 31 vss nmos_5p0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=23090 $Y=1240 $D=2
M11 vss 20 33 vss nmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=24210 $Y=1240 $D=2
M12 20 31 vss vss nmos_5p0 L=6e-07 W=6.23e-06 AD=1.78e-12 AS=1.78e-12 PD=1.112e-05 PS=1.112e-05 NRD=2.24719 NRS=2.24719 m=1 nf=7 $X=26535 $Y=1905 $D=2
M13 vdd wen 29 vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=2545 $Y=4215 $D=8
M14 32 clk vdd vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=3665 $Y=4215 $D=8
M15 2 32 vdd vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=5905 $Y=4215 $D=8
M16 12 wen vdd vdd pmos_5p0 L=6e-07 W=1.488e-05 AD=3.8688e-12 AS=4.7616e-12 PD=1.8e-05 PS=2.368e-05 NRD=0.629032 NRS=0.774194 m=1 nf=6 $X=1260 $Y=9420 $D=8
M17 30 2 29 vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=1.17422e-12 AS=9.988e-13 PD=4.793e-06 PS=5.42e-06 NRD=0.227875 NRS=0.193833 m=1 nf=1 $X=8440 $Y=4215 $D=8
M18 34 32 30 vdd pmos_5p0 L=6e-07 W=9.6e-07 AD=-6.91897e-13 AS=-6.43897e-13 PD=-2.79573e-06 PS=-2.69573e-06 NRD=-0.750757 NRS=-0.698673 m=1 nf=1 $X=10180 $Y=4215 $D=8
M19 vdd 35 34 vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=1.14048e-12 PD=5.42e-06 PS=4.72272e-06 NRD=0.193833 NRS=0.221328 m=1 nf=1 $X=11870 $Y=4215 $D=8
M20 vdd 30 35 vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=14110 $Y=4215 $D=8
M21 16 35 vdd vdd pmos_5p0 L=6e-07 W=5.68e-06 AD=1.4768e-12 AS=2.4992e-12 PD=6.72e-06 PS=1.312e-05 NRD=0.183099 NRS=0.309859 m=1 nf=2 $X=16465 $Y=4215 $D=8
M22 16 32 31 vdd pmos_5p0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=2.13253e-12 PD=5.58e-06 PS=1.01287e-05 NRD=0.229075 NRS=0.413851 m=1 nf=2 $X=19750 $Y=4215 $D=8
M23 33 2 31 vdd pmos_5p0 L=6e-07 W=9.6e-07 AD=-6.59976e-13 AS=-6.40776e-13 PD=-2.72923e-06 PS=-2.68923e-06 NRD=-0.71612 NRS=-0.695287 m=1 nf=1 $X=22550 $Y=5525 $D=8
M24 vdd 20 33 vdd pmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=1.12024e-12 PD=5.42e-06 PS=4.68056e-06 NRD=0.193833 NRS=0.2174 m=1 nf=1 $X=24210 $Y=4215 $D=8
M25 20 31 vdd vdd pmos_5p0 L=6e-07 W=1.54e-05 AD=4.4e-12 AS=4.4e-12 PD=2.16e-05 PS=2.16e-05 NRD=0.909091 NRS=0.909091 m=1 nf=7 $X=26535 $Y=4215 $D=8
X48 vss IGWEN 12 nmos_5p0_CDNS_4025412369678 $T=10115 16070 0 0 $X=9435 $Y=15450
X49 vss GWE 20 nmos_5p0_CDNS_4025412369678 $T=23345 16070 0 0 $X=22665 $Y=15450
X50 vdd IGWEN 12 pmos_5p0_CDNS_4025412369680 $T=10115 9420 0 0 $X=9075 $Y=8800
X51 vdd GWE 20 pmos_5p0_CDNS_4025412369680 $T=23345 9420 0 0 $X=22305 $Y=8800
.ENDS
***************************************
.SUBCKT M1_PACTIVE_CDNS_4025412369650
** N=38 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nmos_1p2$$47641644
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_5p0_CDNS_4025412369671
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT xpredec0_xa 2 3 13 29 30
** N=40 EP=5 IP=40 FDC=4
*.SEEDPROM
M0 40 29 2 3 nmos_5p0 L=6e-07 W=1.225e-05 AD=3.185e-12 AS=7.2275e-12 PD=1.277e-05 PS=2.568e-05 NRD=0.0212245 NRS=0.0481633 m=1 nf=1 $X=3255 $Y=2430 $D=2
M1 3 30 40 3 nmos_5p0 L=6e-07 W=1.225e-05 AD=7.28875e-12 AS=3.185e-12 PD=2.569e-05 PS=1.277e-05 NRD=0.0485714 NRS=0.0212245 m=1 nf=1 $X=4375 $Y=2430 $D=2
M2 2 29 13 13 pmos_5p0 L=6e-07 W=1.52e-05 AD=3.952e-12 AS=6.688e-12 PD=1.572e-05 PS=3.128e-05 NRD=0.0171053 NRS=0.0289474 m=1 nf=1 $X=3255 $Y=19540 $D=8
M3 13 30 2 13 pmos_5p0 L=6e-07 W=1.52e-05 AD=6.688e-12 AS=3.952e-12 PD=3.128e-05 PS=1.572e-05 NRD=0.0289474 NRS=0.0171053 m=1 nf=1 $X=4375 $Y=19540 $D=8
.ENDS
***************************************
.SUBCKT xpredec0_bot 1 2 3 8 9 10 11
** N=33 EP=7 IP=7 FDC=12
M0 2 33 1 1 nmos_5p0 L=6e-07 W=7.04e-06 AD=3.0976e-12 AS=3.0976e-12 PD=1.496e-05 PS=1.496e-05 NRD=0.0625 NRS=0.0625 m=1 nf=1 $X=3755 $Y=35615 $D=2
M1 3 2 1 1 nmos_5p0 L=6e-07 W=5.22e-06 AD=2.2968e-12 AS=2.2968e-12 PD=1.132e-05 PS=1.132e-05 NRD=0.0842912 NRS=0.0842912 m=1 nf=1 $X=6325 $Y=36010 $D=2
M2 2 33 8 8 pmos_5p0 L=6e-07 W=1.769e-05 AD=7.7836e-12 AS=7.7836e-12 PD=3.626e-05 PS=3.626e-05 NRD=0.0248728 NRS=0.0248728 m=1 nf=1 $X=3755 $Y=16320 $D=8
M3 3 2 8 8 pmos_5p0 L=6e-07 W=1.316e-05 AD=5.7904e-12 AS=5.7904e-12 PD=2.72e-05 PS=2.72e-05 NRD=0.0334347 NRS=0.0334347 m=1 nf=1 $X=6325 $Y=20855 $D=8
X4 1 33 9 8 11 10 alatch $T=350 -3160 0 0 $X=-100 $Y=-3165
.ENDS
***************************************
.SUBCKT xpredec0 vss vdd men clk A[1] A[0] x[3] x[2] x[1] x[0]
** N=99 EP=10 IP=158 FDC=56
M0 x[3] 90 vss vss nmos_5p0 L=6e-07 W=1.816e-05 AD=4.7216e-12 AS=5.5388e-12 PD=2.024e-05 PS=2.514e-05 NRD=0.229075 NRS=0.268722 m=1 nf=4 $X=260 $Y=50820 $D=2
M1 x[2] 92 vss vss nmos_5p0 L=6e-07 W=1.816e-05 AD=4.7216e-12 AS=4.7216e-12 PD=2.024e-05 PS=2.024e-05 NRD=0.229075 NRS=0.229075 m=1 nf=4 $X=4740 $Y=50820 $D=2
M2 x[1] 94 vss vss nmos_5p0 L=6e-07 W=1.816e-05 AD=4.7216e-12 AS=4.7216e-12 PD=2.024e-05 PS=2.024e-05 NRD=0.229075 NRS=0.229075 m=1 nf=4 $X=9220 $Y=50820 $D=2
M3 x[0] 96 vss vss nmos_5p0 L=6e-07 W=1.816e-05 AD=4.7216e-12 AS=5.5388e-12 PD=2.024e-05 PS=2.514e-05 NRD=0.229075 NRS=0.268722 m=1 nf=4 $X=13700 $Y=50820 $D=2
M4 17 men vss vss nmos_5p0 L=6e-07 W=1.37e-06 AD=3.562e-13 AS=6.028e-13 PD=1.89e-06 PS=3.62e-06 NRD=0.189781 NRS=0.321168 m=1 nf=1 $X=21630 $Y=51200 $D=2
M5 vss clk 17 vss nmos_5p0 L=6e-07 W=1.37e-06 AD=6.028e-13 AS=3.562e-13 PD=3.62e-06 PS=1.89e-06 NRD=0.321168 NRS=0.189781 m=1 nf=1 $X=22750 $Y=51200 $D=2
M6 x[3] 90 vdd vdd pmos_5p0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.38348e-11 PD=4.744e-05 PS=5.914e-05 NRD=0.0917108 NRS=0.107584 m=1 nf=4 $X=260 $Y=38080 $D=8
M7 x[2] 92 vdd vdd pmos_5p0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.744e-05 PS=4.744e-05 NRD=0.0917108 NRS=0.0917108 m=1 nf=4 $X=4740 $Y=38080 $D=8
M8 x[1] 94 vdd vdd pmos_5p0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.744e-05 PS=4.744e-05 NRD=0.0917108 NRS=0.0917108 m=1 nf=4 $X=9220 $Y=38080 $D=8
M9 x[0] 96 vdd vdd pmos_5p0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.38348e-11 PD=4.744e-05 PS=5.914e-05 NRD=0.0917108 NRS=0.107584 m=1 nf=4 $X=13700 $Y=38080 $D=8
M10 98 men vdd vdd pmos_5p0 L=6e-07 W=1.705e-06 AD=4.39037e-13 AS=1.01447e-12 PD=2.22e-06 PS=4.6e-06 NRD=0.151026 NRS=0.348974 m=1 nf=1 $X=21630 $Y=47525 $D=8
M11 17 clk 98 vdd pmos_5p0 L=6e-07 W=1.705e-06 AD=8.525e-15 AS=-8.525e-15 PD=1e-08 PS=-1e-08 NRD=0.00293255 NRS=-0.00293255 m=1 nf=1 $X=22745 $Y=47525 $D=8
M12 99 clk 17 vdd pmos_5p0 L=6e-07 W=1.705e-06 AD=-8.525e-15 AS=8.525e-15 PD=-1e-08 PS=1e-08 NRD=-0.00293255 NRS=0.00293255 m=1 nf=1 $X=23870 $Y=47525 $D=8
M13 vdd men 99 vdd pmos_5p0 L=6e-07 W=1.705e-06 AD=1.01447e-12 AS=4.39037e-13 PD=4.6e-06 PS=2.22e-06 NRD=0.348974 NRS=0.151026 m=1 nf=1 $X=24985 $Y=47525 $D=8
M14 18 17 vdd vdd pmos_5p0 L=6e-07 W=2.28e-06 AD=5.928e-13 AS=1.0032e-12 PD=3.32e-06 PS=6.32e-06 NRD=0.45614 NRS=0.77193 m=1 nf=2 $X=29010 $Y=47595 $D=8
X17 18 vss 17 vss nmos_1p2$$46563372 $T=29755 51180 0 0 $X=28610 $Y=50495
X18 90 vss vdd 30 31 xpredec0_xa $T=-2205 170 0 0 $X=-1440 $Y=-5
X19 92 vss vdd 30 32 xpredec0_xa $T=11165 170 1 180 $X=3000 $Y=-5
X20 94 vss vdd 33 31 xpredec0_xa $T=6755 170 0 0 $X=7520 $Y=-5
X21 96 vss vdd 33 32 xpredec0_xa $T=20125 170 1 180 $X=11960 $Y=-5
X22 vss 30 33 vdd A[1] 17 18 xpredec0_bot $T=18665 3160 0 0 $X=18135 $Y=-5
X23 vss 31 32 vdd A[0] 17 18 xpredec0_bot $T=27120 3160 0 0 $X=26590 $Y=-5
.ENDS
***************************************
.SUBCKT pmos_5p0_CDNS_4025412369659
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_4025412369658
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ypredec1_ys
** N=8 EP=0 IP=36 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_20 1 2 4 5 7 8
** N=8 EP=6 IP=10 FDC=4
*.SEEDPROM
M0 1 7 4 1 nmos_5p0 L=6e-07 W=2.724e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=3510 $Y=1700 $D=2
M1 8 5 1 1 nmos_5p0 L=6e-07 W=9.08e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=6870 $Y=1700 $D=2
M2 2 7 4 2 pmos_5p0 L=6e-07 W=6e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=3510 $Y=14855 $D=8
M3 8 5 2 2 pmos_5p0 L=6e-07 W=2e-05 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=6870 $Y=14855 $D=8
.ENDS
***************************************
.SUBCKT ICV_21 1 2 4 5 6 7 8 9 11 13
** N=14 EP=10 IP=16 FDC=12
*.SEEDPROM
M0 1 14 6 1 nmos_5p0 L=6e-07 W=2.724e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=9110 $Y=1700 $D=2
M1 12 7 1 1 nmos_5p0 L=6e-07 W=9.08e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=12470 $Y=1700 $D=2
M2 2 14 6 2 pmos_5p0 L=6e-07 W=6e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=9110 $Y=14855 $D=8
M3 12 7 2 2 pmos_5p0 L=6e-07 W=2e-05 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=12470 $Y=14855 $D=8
X4 1 2 4 5 11 14 ICV_20 $T=0 0 0 0 $X=-5 $Y=-5
X5 1 2 8 9 12 13 ICV_20 $T=11200 0 0 0 $X=11195 $Y=-5
.ENDS
***************************************
.SUBCKT pmos_1p2$$47821868
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$47820844
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ypredec1_xa
** N=29 EP=0 IP=36 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_22 1 2 5 8 9 10 11 12
** N=22 EP=8 IP=36 FDC=16
M0 20 10 13 1 nmos_5p0 L=6e-07 W=6.81e-06 AD=1.73655e-12 AS=4.05195e-12 PD=7.32e-06 PS=1.481e-05 NRD=0.0374449 NRS=0.0873715 m=1 nf=1 $X=-2370 $Y=-33035 $D=2
M1 19 9 20 1 nmos_5p0 L=6e-07 W=6.81e-06 AD=3.405e-14 AS=-3.405e-14 PD=1e-08 PS=-1e-08 NRD=0.000734214 NRS=-0.000734214 m=1 nf=1 $X=-1260 $Y=-33035 $D=2
M2 1 2 19 1 nmos_5p0 L=6e-07 W=6.81e-06 AD=3.405e-14 AS=-3.405e-14 PD=1e-08 PS=-1e-08 NRD=0.000734214 NRS=-0.000734214 m=1 nf=1 $X=-140 $Y=-33035 $D=2
M3 1 13 11 1 nmos_5p0 L=6e-07 W=6.81e-06 AD=1.7706e-12 AS=2.1792e-12 PD=8.37e-06 PS=1.1e-05 NRD=0.343612 NRS=0.422907 m=1 nf=3 $X=-2375 $Y=-2950 $D=2
M4 21 5 1 1 nmos_5p0 L=6e-07 W=6.81e-06 AD=-3.405e-14 AS=3.405e-14 PD=-1e-08 PS=1e-08 NRD=-0.000734214 NRS=0.000734214 m=1 nf=1 $X=990 $Y=-33035 $D=2
M5 22 9 21 1 nmos_5p0 L=6e-07 W=6.81e-06 AD=-3.405e-14 AS=3.405e-14 PD=-1e-08 PS=1e-08 NRD=-0.000734214 NRS=0.000734214 m=1 nf=1 $X=2110 $Y=-33035 $D=2
M6 16 10 22 1 nmos_5p0 L=6e-07 W=6.81e-06 AD=4.05195e-12 AS=1.73655e-12 PD=1.481e-05 PS=7.32e-06 NRD=0.0873715 NRS=0.0374449 m=1 nf=1 $X=3220 $Y=-33035 $D=2
M7 12 16 1 1 nmos_5p0 L=6e-07 W=6.81e-06 AD=2.1792e-12 AS=1.7706e-12 PD=1.1e-05 PS=8.37e-06 NRD=0.422907 NRS=0.343612 m=1 nf=3 $X=985 $Y=-2950 $D=2
M8 8 10 13 8 pmos_5p0 L=6e-07 W=5.67e-06 AD=1.4742e-12 AS=2.4948e-12 PD=6.19e-06 PS=1.222e-05 NRD=0.0458554 NRS=0.0776014 m=1 nf=1 $X=-2375 $Y=-19360 $D=8
M9 13 9 8 8 pmos_5p0 L=6e-07 W=5.67e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=-1255 $Y=-19360 $D=8
M10 8 2 13 8 pmos_5p0 L=6e-07 W=5.67e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=-135 $Y=-19360 $D=8
M11 8 13 11 8 pmos_5p0 L=6e-07 W=1.731e-05 AD=4.5006e-12 AS=5.5392e-12 PD=1.887e-05 PS=2.5e-05 NRD=0.135182 NRS=0.166378 m=1 nf=3 $X=-2375 $Y=-10125 $D=8
M12 16 5 8 8 pmos_5p0 L=6e-07 W=5.67e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=985 $Y=-19360 $D=8
M13 8 9 16 8 pmos_5p0 L=6e-07 W=5.67e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=2105 $Y=-19360 $D=8
M14 16 10 8 8 pmos_5p0 L=6e-07 W=5.67e-06 AD=2.4948e-12 AS=1.4742e-12 PD=1.222e-05 PS=6.19e-06 NRD=0.0776014 NRS=0.0458554 m=1 nf=1 $X=3225 $Y=-19360 $D=8
M15 12 16 8 8 pmos_5p0 L=6e-07 W=1.731e-05 AD=5.5392e-12 AS=4.5006e-12 PD=2.5e-05 PS=1.887e-05 NRD=0.166378 NRS=0.135182 m=1 nf=3 $X=985 $Y=-10125 $D=8
.ENDS
***************************************
.SUBCKT ypredec1_bot 1 2 3 10 11 12 13
** N=34 EP=7 IP=20 FDC=12
M0 2 30 1 1 nmos_5p0 L=6e-07 W=4.54e-06 AD=1.9976e-12 AS=1.9976e-12 PD=9.96e-06 PS=9.96e-06 NRD=0.0969163 NRS=0.0969163 m=1 nf=1 $X=3755 $Y=33350 $D=2
M1 3 2 1 1 nmos_5p0 L=6e-07 W=4.54e-06 AD=1.9976e-12 AS=1.9976e-12 PD=9.96e-06 PS=9.96e-06 NRD=0.0969163 NRS=0.0969163 m=1 nf=1 $X=6325 $Y=33350 $D=2
X2 10 2 30 pmos_1p2$$46887980 $T=3910 18340 0 0 $X=2480 $Y=17630
X3 10 3 2 pmos_1p2$$46887980 $T=6480 18340 0 0 $X=5050 $Y=17630
X6 1 30 11 10 13 12 alatch $T=350 -3160 0 0 $X=-100 $Y=-3165
.ENDS
***************************************
.SUBCKT ypredec1 1 2 men clk ly[6] ly[7] ly[0] ly[1] ly[2] ly[3] ly[4] ly[5] ry[0] ry[1] ry[2] ry[3] ry[4] ry[5] ry[6] ry[7]
+ A[2] A[1] A[0]
** N=374 EP=23 IP=151 FDC=172
M0 367 358 1 1 nmos_5p0 L=6e-07 W=9.08e-06 AD=3.9952e-12 AS=3.9952e-12 PD=1.904e-05 PS=1.904e-05 NRD=0.0484581 NRS=0.0484581 m=1 nf=1 $X=2545 $Y=46970 $D=2
M1 1 371 ly[3] 1 nmos_5p0 L=6e-07 W=2.724e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=21585 $Y=46970 $D=2
M2 368 361 1 1 nmos_5p0 L=6e-07 W=9.08e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=24945 $Y=46970 $D=2
M3 188 189 1 1 nmos_5p0 L=6e-07 W=1.36e-06 AD=5.984e-13 AS=5.984e-13 PD=3.6e-06 PS=3.6e-06 NRD=0.323529 NRS=0.323529 m=1 nf=1 $X=31760 $Y=4985 $D=2
M4 189 clk 1 1 nmos_5p0 L=6e-07 W=1.91e-06 AD=4.966e-13 AS=8.404e-13 PD=2.43e-06 PS=4.7e-06 NRD=0.136126 NRS=0.230366 m=1 nf=1 $X=38610 $Y=5010 $D=2
M5 1 men 189 1 nmos_5p0 L=6e-07 W=1.91e-06 AD=8.404e-13 AS=4.966e-13 PD=4.7e-06 PS=2.43e-06 NRD=0.230366 NRS=0.136126 m=1 nf=1 $X=39730 $Y=5010 $D=2
M6 1 372 ly[7] 1 nmos_5p0 L=6e-07 W=2.724e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=43985 $Y=46970 $D=2
M7 369 358 1 1 nmos_5p0 L=6e-07 W=9.08e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=47345 $Y=46970 $D=2
M8 1 373 ry[3] 1 nmos_5p0 L=6e-07 W=2.724e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=66385 $Y=46970 $D=2
M9 370 361 1 1 nmos_5p0 L=6e-07 W=9.08e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=69745 $Y=46970 $D=2
M10 1 374 ry[7] 1 nmos_5p0 L=6e-07 W=2.724e-05 AD=8.7168e-12 AS=8.7168e-12 PD=3.824e-05 PS=3.824e-05 NRD=0.105727 NRS=0.105727 m=1 nf=3 $X=88785 $Y=46970 $D=2
M11 367 358 2 2 pmos_5p0 L=6e-07 W=2e-05 AD=8.8e-12 AS=8.8e-12 PD=4.088e-05 PS=4.088e-05 NRD=0.022 NRS=0.022 m=1 nf=1 $X=2545 $Y=60125 $D=8
M12 2 371 ly[3] 2 pmos_5p0 L=6e-07 W=6e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=21585 $Y=60125 $D=8
M13 368 361 2 2 pmos_5p0 L=6e-07 W=2e-05 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=24945 $Y=60125 $D=8
M14 365 men 2 2 pmos_5p0 L=6e-07 W=2.275e-06 AD=5.915e-13 AS=1.35362e-12 PD=2.795e-06 PS=5.74e-06 NRD=0.114286 NRS=0.261538 m=1 nf=1 $X=36375 $Y=1335 $D=8
M15 189 clk 365 2 pmos_5p0 L=6e-07 W=2.275e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=37495 $Y=1335 $D=8
M16 366 clk 189 2 pmos_5p0 L=6e-07 W=2.275e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=38615 $Y=1335 $D=8
M17 2 men 366 2 pmos_5p0 L=6e-07 W=2.275e-06 AD=1.34225e-12 AS=5.915e-13 PD=5.73e-06 PS=2.795e-06 NRD=0.259341 NRS=0.114286 m=1 nf=1 $X=39735 $Y=1335 $D=8
M18 2 372 ly[7] 2 pmos_5p0 L=6e-07 W=6e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=43985 $Y=60125 $D=8
M19 369 358 2 2 pmos_5p0 L=6e-07 W=2e-05 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=47345 $Y=60125 $D=8
M20 2 373 ry[3] 2 pmos_5p0 L=6e-07 W=6e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=66385 $Y=60125 $D=8
M21 370 361 2 2 pmos_5p0 L=6e-07 W=2e-05 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=69745 $Y=60125 $D=8
M22 2 374 ry[7] 2 pmos_5p0 L=6e-07 W=6e-05 AD=1.92e-11 AS=1.92e-11 PD=8.192e-05 PS=8.192e-05 NRD=0.048 NRS=0.048 m=1 nf=3 $X=88785 $Y=60125 $D=8
X26 2 188 189 pmos_1p2$$47109164 $T=32795 1405 1 180 $X=28795 $Y=720
X27 1 2 ly[0] 357 ly[1] 359 ly[2] 360 367 371 ICV_21 $T=1275 45270 0 0 $X=1270 $Y=45265
X28 1 2 ly[4] 362 ly[5] 363 ly[6] 364 368 372 ICV_21 $T=23675 45270 0 0 $X=23670 $Y=45265
X29 1 2 ry[0] 357 ry[1] 359 ry[2] 360 369 373 ICV_21 $T=46075 45270 0 0 $X=46070 $Y=45265
X30 1 2 ry[4] 362 ry[5] 363 ry[6] 364 370 374 ICV_21 $T=68475 45270 0 0 $X=68470 $Y=45265
X31 1 195 194 2 192 190 363 364 ICV_22 $T=33645 42985 1 180 $X=28115 $Y=7365
X32 1 195 194 2 193 190 361 362 ICV_22 $T=41810 42985 1 180 $X=36280 $Y=7365
X33 1 195 194 2 192 191 359 360 ICV_22 $T=49980 42985 1 180 $X=44450 $Y=7365
X34 1 195 194 2 193 191 358 357 ICV_22 $T=58150 42985 1 180 $X=52620 $Y=7365
X35 1 190 191 2 A[2] 189 188 ypredec1_bot $T=1920 5135 0 0 $X=1820 $Y=1970
X36 1 192 193 2 A[1] 189 188 ypredec1_bot $T=10375 5135 0 0 $X=10275 $Y=1970
X37 1 194 195 2 A[0] 189 188 ypredec1_bot $T=18830 5135 0 0 $X=18730 $Y=1970
.ENDS
***************************************
.SUBCKT M1_PSUB_CDNS_4025412369616
** N=2401 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pmoscap_W2_5_R270
** N=13 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmoscap_W2_5_477_R270
** N=26 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_23
** N=6 EP=0 IP=8 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT M1_NWELL$$204218412
** N=49 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_PACTIVE$$204148780
** N=13 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_40254123696102 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 2 nmos_5p0 L=6e-07 W=1.011e-05 AD=4.4484e-12 AS=4.4484e-12 PD=2.11e-05 PS=2.11e-05 NRD=0.0435213 NRS=0.0435213 m=1 nf=1 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT pmos_1p2$$204216364_R90 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pmos_5p0 L=6e-07 W=2.526e-05 AD=6.5676e-12 AS=1.11144e-11 PD=2.63e-05 PS=5.228e-05 NRD=0.0411718 NRS=0.0696754 m=1 nf=2 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT pmos_5p0_CDNS_40254123696100 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 pmos_5p0 L=6e-07 W=6.59e-06 AD=2.8996e-12 AS=2.8996e-12 PD=1.406e-05 PS=1.406e-05 NRD=0.0667678 NRS=0.0667678 m=1 nf=1 $X=0 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_40254123696111 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 2 nmos_5p0 L=6e-07 W=2.64e-06 AD=1.1616e-12 AS=1.1616e-12 PD=6.16e-06 PS=6.16e-06 NRD=0.166667 NRS=0.166667 m=1 nf=1 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT pmos_5p0_CDNS_40254123696105
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT M1_POLY2_CDNS_40254123696102
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nmos_5p0_CDNS_40254123696108
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$49272876_R270 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pmos_5p0 L=6e-07 W=1.1e-05 AD=2.86e-12 AS=4.84e-12 PD=1.204e-05 PS=2.376e-05 NRD=0.0945455 NRS=0.16 m=1 nf=2 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT pmos_5p0_CDNS_40254123696106
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT xdec 1 2 men 6 vss 8 28 vdd
** N=98 EP=8 IP=41 FDC=6
*.SEEDPROM
M0 2 6 men vss nmos_5p0 L=6e-07 W=6.6e-06 AD=2.904e-12 AS=1.716e-12 PD=1.496e-05 PS=7.64e-06 NRD=0.266667 NRS=0.157576 m=1 nf=2 $X=37460 $Y=965 $D=2
M1 vss 8 6 vss nmos_5p0 L=6e-07 W=6.6e-07 AD=2.904e-13 AS=2.904e-13 PD=2.2e-06 PS=2.2e-06 NRD=0.666667 NRS=0.666667 m=1 nf=1 $X=45970 $Y=965 $D=2
M2 2 8 men vdd pmos_5p0 L=6e-07 W=6.6e-06 AD=2.904e-12 AS=1.716e-12 PD=1.496e-05 PS=7.64e-06 NRD=0.266667 NRS=0.157576 m=1 nf=2 $X=32185 $Y=965 $D=8
M3 vdd 8 6 vdd pmos_5p0 L=6e-07 W=1.59e-06 AD=6.996e-13 AS=6.996e-13 PD=4.06e-06 PS=4.06e-06 NRD=0.27673 NRS=0.27673 m=1 nf=1 $X=43020 $Y=965 $D=8
X12 vdd 1 2 pmos_1p2$$49272876_R270 $T=29780 1120 0 90 $X=23605 $Y=-360
X13 vdd 28 2 pmos_1p2$$49272876_R270 $T=91805 1120 1 90 $X=91120 $Y=-360
.ENDS
***************************************
.SUBCKT ICV_24 1 50 94 95 96 100 101 114 117 118 121
** N=125 EP=11 IP=142 FDC=12
*.SEEDPROM
X0 114 94 95 115 1 96 117 50 xdec $T=0 0 1 0 $X=-5 $Y=-5640
X1 118 100 95 119 1 101 121 50 xdec $T=0 0 0 0 $X=-5 $Y=-1115
.ENDS
***************************************
.SUBCKT xdec8_64 men vss DRWL vdd xa[0] xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] xa[7] LWL[0] LWL[1] LWL[2] LWL[3] LWL[4] LWL[5] LWL[6] LWL[7]
+ RWL[1] RWL[2] RWL[4] RWL[6] RWL[7] RWL[3] RWL[5] RWL[0]
** N=317 EP=28 IP=541 FDC=156
M0 vss 288 LWL[0] vss nmos_5p0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=24970 $Y=260 $D=2
M1 288 272 vss vss nmos_5p0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=24970 $Y=2660 $D=2
M2 vss 270 286 vss nmos_5p0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=24970 $Y=5740 $D=2
M3 vss 286 LWL[1] vss nmos_5p0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=24970 $Y=7020 $D=2
M4 vss 292 LWL[2] vss nmos_5p0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=24970 $Y=9260 $D=2
M5 292 276 vss vss nmos_5p0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=24970 $Y=11660 $D=2
M6 vss 274 290 vss nmos_5p0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=24970 $Y=14740 $D=2
M7 vss 290 LWL[3] vss nmos_5p0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=24970 $Y=16020 $D=2
M8 vss 296 LWL[4] vss nmos_5p0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=24970 $Y=18260 $D=2
M9 296 280 vss vss nmos_5p0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=24970 $Y=20660 $D=2
M10 vss 278 294 vss nmos_5p0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=24970 $Y=23740 $D=2
M11 vss 294 LWL[5] vss nmos_5p0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=24970 $Y=25020 $D=2
M12 vss 300 LWL[6] vss nmos_5p0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=24970 $Y=27260 $D=2
M13 300 284 vss vss nmos_5p0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=24970 $Y=29660 $D=2
M14 vss 282 298 vss nmos_5p0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=24970 $Y=32740 $D=2
M15 vss 298 LWL[7] vss nmos_5p0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=24970 $Y=34020 $D=2
M16 272 273 vss vss nmos_5p0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=9.68e-13 PD=5.28e-06 PS=5.28e-06 NRD=0.2 NRS=0.2 m=1 nf=1 $X=55250 $Y=260 $D=2
M17 vss 271 270 vss nmos_5p0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=55250 $Y=8140 $D=2
M18 276 277 vss vss nmos_5p0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=55250 $Y=9260 $D=2
M19 vss 275 274 vss nmos_5p0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=55250 $Y=17140 $D=2
M20 280 281 vss vss nmos_5p0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=55250 $Y=18260 $D=2
M21 vss 279 278 vss nmos_5p0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=55250 $Y=26140 $D=2
M22 284 285 vss vss nmos_5p0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=55250 $Y=27260 $D=2
M23 vss 283 282 vss nmos_5p0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=9.68e-13 PD=5.28e-06 PS=5.28e-06 NRD=0.2 NRS=0.2 m=1 nf=1 $X=55250 $Y=35140 $D=2
M24 29 vdd men vss nmos_5p0 L=6e-07 W=6.59e-06 AD=2.8996e-12 AS=2.8996e-12 PD=1.406e-05 PS=1.406e-05 NRD=0.0667678 NRS=0.0667678 m=1 nf=1 $X=61430 $Y=38365 $D=2
M25 305 vdd vss vss nmos_5p0 L=6e-07 W=3.15e-06 AD=7.32375e-13 AS=2.079e-12 PD=3.615e-06 PS=7.62e-06 NRD=0.0738095 NRS=0.209524 m=1 nf=1 $X=75090 $Y=315 $D=2
M26 304 vdd 305 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=75090 $Y=1380 $D=2
M27 273 xa[0] 304 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=75090 $Y=2500 $D=2
M28 302 xa[1] 271 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=75090 $Y=5900 $D=2
M29 303 vdd 302 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=75090 $Y=7020 $D=2
M30 vss vdd 303 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=75090 $Y=8085 $D=2
M31 309 vdd vss vss nmos_5p0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=75090 $Y=9315 $D=2
M32 308 vdd 309 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=75090 $Y=10380 $D=2
M33 277 xa[2] 308 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=75090 $Y=11500 $D=2
M34 306 xa[3] 275 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=75090 $Y=14900 $D=2
M35 307 vdd 306 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=75090 $Y=16020 $D=2
M36 vss vdd 307 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=75090 $Y=17085 $D=2
M37 313 vdd vss vss nmos_5p0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=75090 $Y=18315 $D=2
M38 312 vdd 313 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=75090 $Y=19380 $D=2
M39 281 xa[4] 312 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=75090 $Y=20500 $D=2
M40 310 xa[5] 279 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=75090 $Y=23900 $D=2
M41 311 vdd 310 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=75090 $Y=25020 $D=2
M42 vss vdd 311 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=75090 $Y=26085 $D=2
M43 317 vdd vss vss nmos_5p0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=75090 $Y=27315 $D=2
M44 316 vdd 317 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=75090 $Y=28380 $D=2
M45 285 xa[6] 316 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=75090 $Y=29500 $D=2
M46 314 xa[7] 283 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=75090 $Y=32900 $D=2
M47 315 vdd 314 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=75090 $Y=34020 $D=2
M48 vss vdd 315 vss nmos_5p0 L=6e-07 W=3.15e-06 AD=2.079e-12 AS=7.32375e-13 PD=7.62e-06 PS=3.615e-06 NRD=0.209524 NRS=0.0738095 m=1 nf=1 $X=75090 $Y=35085 $D=2
M49 vss 289 RWL[0] vss nmos_5p0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=108885 $Y=260 $D=2
M50 289 272 vss vss nmos_5p0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=108885 $Y=2660 $D=2
M51 vss 270 287 vss nmos_5p0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=108885 $Y=5740 $D=2
M52 vss 287 RWL[1] vss nmos_5p0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=108885 $Y=7020 $D=2
M53 vss 293 RWL[2] vss nmos_5p0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=108885 $Y=9260 $D=2
M54 293 276 vss vss nmos_5p0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=108885 $Y=11660 $D=2
M55 vss 274 291 vss nmos_5p0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=108885 $Y=14740 $D=2
M56 vss 291 RWL[3] vss nmos_5p0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=108885 $Y=16020 $D=2
M57 vss 297 RWL[4] vss nmos_5p0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=108885 $Y=18260 $D=2
M58 297 280 vss vss nmos_5p0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=108885 $Y=20660 $D=2
M59 vss 278 295 vss nmos_5p0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=108885 $Y=23740 $D=2
M60 vss 295 RWL[5] vss nmos_5p0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=108885 $Y=25020 $D=2
M61 vss 301 RWL[6] vss nmos_5p0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=108885 $Y=27260 $D=2
M62 301 284 vss vss nmos_5p0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=108885 $Y=29660 $D=2
M63 vss 282 299 vss nmos_5p0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=108885 $Y=32740 $D=2
M64 vss 299 RWL[7] vss nmos_5p0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=108885 $Y=34020 $D=2
M65 vdd vss vdd vdd pmos_5p0 L=3.94e-06 W=4.9455e-05 AD=0 AS=3.14863e-11 PD=0 PS=0.00012136 NRD=0 NRS=1.04277 m=1 nf=9 $X=2985 $Y=280 $D=8
M66 vdd 288 LWL[0] vdd pmos_5p0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=13295 $Y=260 $D=8
M67 LWL[1] 286 vdd vdd pmos_5p0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=13295 $Y=5900 $D=8
M68 vdd 292 LWL[2] vdd pmos_5p0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=13295 $Y=9260 $D=8
M69 LWL[3] 290 vdd vdd pmos_5p0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=13295 $Y=14900 $D=8
M70 vdd 296 LWL[4] vdd pmos_5p0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=13295 $Y=18260 $D=8
M71 LWL[5] 294 vdd vdd pmos_5p0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=13295 $Y=23900 $D=8
M72 vdd 300 LWL[6] vdd pmos_5p0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=13295 $Y=27260 $D=8
M73 LWL[7] 298 vdd vdd pmos_5p0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=13295 $Y=32900 $D=8
M74 vdd vdd 273 vdd pmos_5p0 L=6e-07 W=5.24e-06 AD=1.834e-12 AS=1.3624e-12 PD=9.26e-06 PS=6.28e-06 NRD=0.267176 NRS=0.198473 m=1 nf=2 $X=80610 $Y=260 $D=8
M75 273 xa[0] vdd vdd pmos_5p0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=80610 $Y=2500 $D=8
M76 vdd xa[1] 271 vdd pmos_5p0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=80610 $Y=5900 $D=8
M77 vdd vdd 271 vdd pmos_5p0 L=6e-07 W=5.24e-06 AD=1.3624e-12 AS=1.3624e-12 PD=6.28e-06 PS=6.28e-06 NRD=0.198473 NRS=0.198473 m=1 nf=2 $X=80610 $Y=7020 $D=8
M78 vdd vdd 277 vdd pmos_5p0 L=6e-07 W=5.24e-06 AD=1.3624e-12 AS=1.3624e-12 PD=6.28e-06 PS=6.28e-06 NRD=0.198473 NRS=0.198473 m=1 nf=2 $X=80610 $Y=9260 $D=8
M79 277 xa[2] vdd vdd pmos_5p0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=80610 $Y=11500 $D=8
M80 vdd xa[3] 275 vdd pmos_5p0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=80610 $Y=14900 $D=8
M81 vdd vdd 275 vdd pmos_5p0 L=6e-07 W=5.24e-06 AD=1.3624e-12 AS=1.3624e-12 PD=6.28e-06 PS=6.28e-06 NRD=0.198473 NRS=0.198473 m=1 nf=2 $X=80610 $Y=16020 $D=8
M82 vdd vdd 281 vdd pmos_5p0 L=6e-07 W=5.24e-06 AD=1.3624e-12 AS=1.3624e-12 PD=6.28e-06 PS=6.28e-06 NRD=0.198473 NRS=0.198473 m=1 nf=2 $X=80610 $Y=18260 $D=8
M83 281 xa[4] vdd vdd pmos_5p0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=80610 $Y=20500 $D=8
M84 vdd xa[5] 279 vdd pmos_5p0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=80610 $Y=23900 $D=8
M85 vdd vdd 279 vdd pmos_5p0 L=6e-07 W=5.24e-06 AD=1.3624e-12 AS=1.3624e-12 PD=6.28e-06 PS=6.28e-06 NRD=0.198473 NRS=0.198473 m=1 nf=2 $X=80610 $Y=25020 $D=8
M86 vdd vdd 285 vdd pmos_5p0 L=6e-07 W=5.24e-06 AD=1.3624e-12 AS=1.3624e-12 PD=6.28e-06 PS=6.28e-06 NRD=0.198473 NRS=0.198473 m=1 nf=2 $X=80610 $Y=27260 $D=8
M87 285 xa[6] vdd vdd pmos_5p0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=80610 $Y=29500 $D=8
M88 vdd xa[7] 283 vdd pmos_5p0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=80610 $Y=32900 $D=8
M89 vdd vdd 283 vdd pmos_5p0 L=6e-07 W=5.24e-06 AD=1.834e-12 AS=1.3624e-12 PD=9.26e-06 PS=6.28e-06 NRD=0.267176 NRS=0.198473 m=1 nf=2 $X=80610 $Y=34020 $D=8
M90 vdd 289 RWL[0] vdd pmos_5p0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=115560 $Y=260 $D=8
M91 RWL[1] 287 vdd vdd pmos_5p0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=115560 $Y=5900 $D=8
M92 vdd 293 RWL[2] vdd pmos_5p0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=115560 $Y=9260 $D=8
M93 RWL[3] 291 vdd vdd pmos_5p0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=115560 $Y=14900 $D=8
M94 vdd 297 RWL[4] vdd pmos_5p0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=115560 $Y=18260 $D=8
M95 RWL[5] 295 vdd vdd pmos_5p0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=115560 $Y=23900 $D=8
M96 vdd 301 RWL[6] vdd pmos_5p0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=115560 $Y=27260 $D=8
M97 RWL[7] 299 vdd vdd pmos_5p0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=115560 $Y=32900 $D=8
M98 vdd vss vdd vdd pmos_5p0 L=3.94e-06 W=4.9455e-05 AD=0 AS=3.14863e-11 PD=0 PS=0.00012136 NRD=0 NRS=1.04277 m=1 nf=9 $X=130365 $Y=280 $D=8
X110 DLWL vss 37 nmos_5p0_CDNS_40254123696102 $T=31730 38360 0 90 $X=21000 $Y=37680
X111 DRWL vss 38 nmos_5p0_CDNS_40254123696102 $T=116730 38360 0 90 $X=106000 $Y=37680
X112 vdd DLWL 37 pmos_1p2$$204216364_R90 $T=46225 38515 0 90 $X=32935 $Y=37035
X113 vdd DRWL 38 pmos_1p2$$204216364_R90 $T=104750 38515 0 90 $X=91460 $Y=37035
X114 37 vdd 29 vdd pmos_5p0_CDNS_40254123696100 $T=55020 38360 0 90 $X=47810 $Y=37320
X115 men 29 vss vdd pmos_5p0_CDNS_40254123696100 $T=76520 38360 0 90 $X=69310 $Y=37320
X116 38 vdd 29 vdd pmos_5p0_CDNS_40254123696100 $T=89870 38360 0 90 $X=82660 $Y=37320
X117 37 vss 29 nmos_5p0_CDNS_40254123696111 $T=59565 38360 0 90 $X=56305 $Y=37680
X118 38 vss 29 nmos_5p0_CDNS_40254123696111 $T=81415 38360 0 90 $X=78155 $Y=37680
X119 vss vdd 270 men 271 272 273 286 287 288 289 ICV_24 $T=8635 4500 1 0 $X=8630 $Y=-1140
X120 vss vdd 274 men 275 276 277 290 291 292 293 ICV_24 $T=8635 13500 1 0 $X=8630 $Y=7860
X121 vss vdd 278 men 279 280 281 294 295 296 297 ICV_24 $T=8635 22500 1 0 $X=8630 $Y=16860
X122 vss vdd 282 men 283 284 285 298 299 300 301 ICV_24 $T=8635 31500 1 0 $X=8630 $Y=25860
.ENDS
***************************************
.SUBCKT 018SRAM_cell1_cutPC
** N=7 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT 018SRAM_strap1_2x_bndry
** N=13 EP=0 IP=12 FDC=0
.ENDS
***************************************
.SUBCKT ICV_25 1 2 10 13 14 15 16
** N=16 EP=7 IP=27 FDC=8
*.SEEDPROM
M0 2 10 14 10 nmos_5p0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=3180 $Y=-1030 $D=2
M1 16 10 2 10 nmos_5p0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=3180 $Y=260 $D=2
M2 10 13 14 10 nmos_5p0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=3630 $Y=-2660 $D=2
M3 10 15 16 10 nmos_5p0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=3630 $Y=1710 $D=2
M4 13 14 10 10 nmos_5p0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=4770 $Y=-2660 $D=2
M5 15 16 10 10 nmos_5p0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=4770 $Y=1710 $D=2
M6 1 10 13 10 nmos_5p0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=5220 $Y=-1030 $D=2
M7 15 10 1 10 nmos_5p0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=5220 $Y=260 $D=2
.ENDS
***************************************
.SUBCKT ICV_26 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 35 36
+ 37 38 39 40 41 42
** N=66 EP=26 IP=87 FDC=208
*.SEEDPROM
M0 1 22 20 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-8370 $Y=3560 $D=8
M1 1 44 43 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-8370 $Y=4840 $D=8
M2 1 48 47 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-8370 $Y=21560 $D=8
M3 1 60 59 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-8370 $Y=22840 $D=8
M4 22 20 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-7230 $Y=3560 $D=8
M5 44 43 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-7230 $Y=4840 $D=8
M6 48 47 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-7230 $Y=21560 $D=8
M7 60 59 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-7230 $Y=22840 $D=8
M8 1 26 24 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-5370 $Y=3560 $D=8
M9 1 46 45 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-5370 $Y=4840 $D=8
M10 1 50 49 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-5370 $Y=21560 $D=8
M11 1 62 61 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-5370 $Y=22840 $D=8
M12 26 24 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-4230 $Y=3560 $D=8
M13 46 45 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-4230 $Y=4840 $D=8
M14 50 49 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-4230 $Y=21560 $D=8
M15 62 61 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-4230 $Y=22840 $D=8
M16 1 30 28 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=3560 $D=8
M17 1 52 51 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=4840 $D=8
M18 1 56 55 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=21560 $D=8
M19 1 64 63 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=22840 $D=8
M20 30 28 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=3560 $D=8
M21 52 51 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=4840 $D=8
M22 56 55 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=21560 $D=8
M23 64 63 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=22840 $D=8
M24 1 34 32 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=3560 $D=8
M25 1 54 53 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=4840 $D=8
M26 1 58 57 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=21560 $D=8
M27 1 66 65 1 pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=22840 $D=8
M28 34 32 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=3560 $D=8
M29 54 53 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=4840 $D=8
M30 58 57 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=21560 $D=8
M31 66 65 1 1 pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=22840 $D=8
X32 1 2 3 4 5 6 11 12 13 14 15 16 17 18 43 44 45 46 47 48
+ 49 50 51 52 53 54 55 56 57 58
+ ICV_5 $T=0 4500 0 0 $X=-9340 $Y=4160
X33 1 2 7 8 9 10 11 12 13 14 15 16 17 18 59 60 61 62 35 36
+ 37 38 63 64 65 66 39 40 41 42
+ ICV_5 $T=0 22500 0 0 $X=-9340 $Y=22160
X34 2 2 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 ICV_8 $T=0 0 0 0 $X=-9340 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_27
** N=19 EP=0 IP=30 FDC=0
.ENDS
***************************************
.SUBCKT ICV_28
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT lcol4_64 VSS VDD WEN[2] pcb[2] b[23] bb[23] men WEN[0] pcb[0] b[7] bb[7] WEN[3] pcb[3] b[24] bb[24] WEN[1] pcb[1] b[8] bb[8] WL[0]
+ WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] GWEN GWE ypass[0] ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] din[1] q[1] din[3]
+ q[3] din[0] q[0] din[2] q[2] b[26] bb[26] bb[27] b[27] bb[25] b[25] b[10] bb[10] bb[11] b[11] bb[9] b[9] b[28] bb[28] bb[29]
+ b[29] b[30] bb[30] bb[31] b[31] b[20] bb[20] bb[21] b[21] b[22] bb[22] b[16] bb[16] bb[17] b[17] b[18] bb[18] bb[19] b[19] b[12]
+ bb[12] bb[13] b[13] b[14] bb[14] bb[15] b[15] b[0] bb[0] bb[1] b[1] b[2] bb[2] bb[3] b[3] b[4] bb[4] bb[5] b[5] b[6]
+ bb[6]
** N=500 EP=101 IP=1003 FDC=2761
*.SEEDPROM
M0 138 VSS 47 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=105785 $Y=151295 $D=2
M1 47 VSS 140 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=105785 $Y=195005 $D=2
M2 VSS 137 138 VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=106235 $Y=152745 $D=2
M3 VSS 139 140 VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=106235 $Y=193375 $D=2
M4 137 138 VSS VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=107375 $Y=152745 $D=2
M5 139 140 VSS VSS nmos_5p0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=107375 $Y=193375 $D=2
M6 137 VSS 46 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=107825 $Y=151295 $D=2
M7 46 VSS 139 VSS nmos_5p0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=107825 $Y=195005 $D=2
M8 VDD 186 188 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-1765 $Y=154595 $D=8
M9 VDD 344 343 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-1765 $Y=155875 $D=8
M10 VDD 352 351 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-1765 $Y=190595 $D=8
M11 VDD 202 204 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-1765 $Y=191875 $D=8
M12 186 188 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-625 $Y=154595 $D=8
M13 344 343 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-625 $Y=155875 $D=8
M14 352 351 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-625 $Y=190595 $D=8
M15 202 204 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-625 $Y=191875 $D=8
M16 439 ypass[7] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=-770 $Y=87735 $D=8
M17 VDD 182 184 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=1235 $Y=154595 $D=8
M18 VDD 346 345 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=1235 $Y=155875 $D=8
M19 VDD 354 353 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=1235 $Y=190595 $D=8
M20 VDD 198 200 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=1235 $Y=191875 $D=8
M21 182 184 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=2375 $Y=154595 $D=8
M22 346 345 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=2375 $Y=155875 $D=8
M23 354 353 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=2375 $Y=190595 $D=8
M24 198 200 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=2375 $Y=191875 $D=8
M25 440 ypass[6] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=1760 $Y=87735 $D=8
M26 VDD 178 180 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=4235 $Y=154595 $D=8
M27 VDD 348 347 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=4235 $Y=155875 $D=8
M28 VDD 356 355 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=4235 $Y=190595 $D=8
M29 VDD 194 196 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=4235 $Y=191875 $D=8
M30 178 180 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=5375 $Y=154595 $D=8
M31 348 347 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=5375 $Y=155875 $D=8
M32 356 355 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=5375 $Y=190595 $D=8
M33 194 196 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=5375 $Y=191875 $D=8
M34 441 ypass[5] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=5425 $Y=87735 $D=8
M35 VDD 174 176 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=7235 $Y=154595 $D=8
M36 VDD 350 349 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=7235 $Y=155875 $D=8
M37 VDD 358 357 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=7235 $Y=190595 $D=8
M38 VDD 190 192 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=7235 $Y=191875 $D=8
M39 174 176 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=8375 $Y=154595 $D=8
M40 350 349 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=8375 $Y=155875 $D=8
M41 358 357 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=8375 $Y=190595 $D=8
M42 190 192 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=8375 $Y=191875 $D=8
M43 442 ypass[4] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=7955 $Y=87735 $D=8
M44 VDD 146 148 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=10235 $Y=154595 $D=8
M45 VDD 360 359 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=10235 $Y=155875 $D=8
M46 VDD 368 367 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=10235 $Y=190595 $D=8
M47 VDD 218 220 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=10235 $Y=191875 $D=8
M48 146 148 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=11375 $Y=154595 $D=8
M49 360 359 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=11375 $Y=155875 $D=8
M50 368 367 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=11375 $Y=190595 $D=8
M51 218 220 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=11375 $Y=191875 $D=8
M52 443 ypass[3] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=11615 $Y=87735 $D=8
M53 VDD 142 144 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=13235 $Y=154595 $D=8
M54 VDD 362 361 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=13235 $Y=155875 $D=8
M55 VDD 370 369 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=13235 $Y=190595 $D=8
M56 VDD 214 216 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=13235 $Y=191875 $D=8
M57 142 144 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=14375 $Y=154595 $D=8
M58 362 361 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=14375 $Y=155875 $D=8
M59 370 369 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=14375 $Y=190595 $D=8
M60 214 216 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=14375 $Y=191875 $D=8
M61 444 ypass[2] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=14145 $Y=87735 $D=8
M62 VDD 154 156 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=16235 $Y=154595 $D=8
M63 VDD 364 363 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=16235 $Y=155875 $D=8
M64 VDD 372 371 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=16235 $Y=190595 $D=8
M65 VDD 210 212 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=16235 $Y=191875 $D=8
M66 154 156 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=17375 $Y=154595 $D=8
M67 364 363 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=17375 $Y=155875 $D=8
M68 372 371 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=17375 $Y=190595 $D=8
M69 210 212 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=17375 $Y=191875 $D=8
M70 445 ypass[1] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=17810 $Y=87735 $D=8
M71 VDD 150 152 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=19235 $Y=154595 $D=8
M72 VDD 366 365 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=19235 $Y=155875 $D=8
M73 VDD 374 373 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=19235 $Y=190595 $D=8
M74 VDD 206 208 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=19235 $Y=191875 $D=8
M75 150 152 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=20375 $Y=154595 $D=8
M76 366 365 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=20375 $Y=155875 $D=8
M77 374 373 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=20375 $Y=190595 $D=8
M78 206 208 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=20375 $Y=191875 $D=8
M79 327 ypass[0] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=20340 $Y=87735 $D=8
M80 VDD 475 476 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=25235 $Y=190595 $D=8
M81 VDD 234 236 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=25235 $Y=191875 $D=8
M82 325 ypass[7] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=24015 $Y=87735 $D=8
M83 475 476 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=26375 $Y=190595 $D=8
M84 234 236 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=26375 $Y=191875 $D=8
M85 335 ypass[6] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=26540 $Y=87735 $D=8
M86 VDD 473 474 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=28235 $Y=190595 $D=8
M87 VDD 230 232 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=28235 $Y=191875 $D=8
M88 473 474 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=29375 $Y=190595 $D=8
M89 230 232 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=29375 $Y=191875 $D=8
M90 VDD 471 472 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=31235 $Y=190595 $D=8
M91 VDD 226 228 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=31235 $Y=191875 $D=8
M92 334 ypass[5] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=30205 $Y=87735 $D=8
M93 471 472 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=32375 $Y=190595 $D=8
M94 226 228 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=32375 $Y=191875 $D=8
M95 333 ypass[4] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=32735 $Y=87735 $D=8
M96 VDD 469 470 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=34235 $Y=190595 $D=8
M97 VDD 222 224 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=34235 $Y=191875 $D=8
M98 469 470 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=35375 $Y=190595 $D=8
M99 222 224 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=35375 $Y=191875 $D=8
M100 VDD 483 484 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=37235 $Y=190595 $D=8
M101 VDD 250 252 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=37235 $Y=191875 $D=8
M102 332 ypass[3] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=36395 $Y=87735 $D=8
M103 483 484 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=38375 $Y=190595 $D=8
M104 250 252 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=38375 $Y=191875 $D=8
M105 331 ypass[2] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=38925 $Y=87735 $D=8
M106 VDD 481 482 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=40235 $Y=190595 $D=8
M107 VDD 246 248 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=40235 $Y=191875 $D=8
M108 481 482 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=41375 $Y=190595 $D=8
M109 246 248 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=41375 $Y=191875 $D=8
M110 VDD 479 480 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=43235 $Y=190595 $D=8
M111 VDD 242 244 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=43235 $Y=191875 $D=8
M112 330 ypass[1] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=42590 $Y=87735 $D=8
M113 479 480 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=44375 $Y=190595 $D=8
M114 242 244 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=44375 $Y=191875 $D=8
M115 VDD 477 478 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=46235 $Y=190595 $D=8
M116 VDD 238 240 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=46235 $Y=191875 $D=8
M117 329 ypass[0] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=45120 $Y=87735 $D=8
M118 477 478 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=47375 $Y=190595 $D=8
M119 238 240 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=47375 $Y=191875 $D=8
M120 VDD 266 268 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=52235 $Y=154595 $D=8
M121 VDD 376 375 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=52235 $Y=155875 $D=8
M122 VDD 384 383 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=52235 $Y=190595 $D=8
M123 VDD 413 414 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=52235 $Y=191875 $D=8
M124 266 268 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=53375 $Y=154595 $D=8
M125 376 375 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=53375 $Y=155875 $D=8
M126 384 383 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=53375 $Y=190595 $D=8
M127 413 414 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=53375 $Y=191875 $D=8
M128 446 ypass[7] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=53230 $Y=87735 $D=8
M129 VDD 262 264 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=55235 $Y=154595 $D=8
M130 VDD 378 377 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=55235 $Y=155875 $D=8
M131 VDD 386 385 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=55235 $Y=190595 $D=8
M132 VDD 411 412 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=55235 $Y=191875 $D=8
M133 262 264 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=56375 $Y=154595 $D=8
M134 378 377 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=56375 $Y=155875 $D=8
M135 386 385 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=56375 $Y=190595 $D=8
M136 411 412 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=56375 $Y=191875 $D=8
M137 447 ypass[6] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=55760 $Y=87735 $D=8
M138 VDD 258 260 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=58235 $Y=154595 $D=8
M139 VDD 380 379 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=58235 $Y=155875 $D=8
M140 VDD 388 387 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=58235 $Y=190595 $D=8
M141 VDD 409 410 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=58235 $Y=191875 $D=8
M142 258 260 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=59375 $Y=154595 $D=8
M143 380 379 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=59375 $Y=155875 $D=8
M144 388 387 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=59375 $Y=190595 $D=8
M145 409 410 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=59375 $Y=191875 $D=8
M146 448 ypass[5] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=59425 $Y=87735 $D=8
M147 VDD 254 256 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=61235 $Y=154595 $D=8
M148 VDD 382 381 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=61235 $Y=155875 $D=8
M149 VDD 390 389 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=61235 $Y=190595 $D=8
M150 VDD 407 408 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=61235 $Y=191875 $D=8
M151 254 256 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=62375 $Y=154595 $D=8
M152 382 381 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=62375 $Y=155875 $D=8
M153 390 389 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=62375 $Y=190595 $D=8
M154 407 408 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=62375 $Y=191875 $D=8
M155 449 ypass[4] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=61955 $Y=87735 $D=8
M156 VDD 162 164 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=64235 $Y=154595 $D=8
M157 VDD 392 391 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=64235 $Y=155875 $D=8
M158 VDD 400 399 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=64235 $Y=190595 $D=8
M159 VDD 421 422 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=64235 $Y=191875 $D=8
M160 162 164 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=65375 $Y=154595 $D=8
M161 392 391 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=65375 $Y=155875 $D=8
M162 400 399 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=65375 $Y=190595 $D=8
M163 421 422 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=65375 $Y=191875 $D=8
M164 450 ypass[3] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=65615 $Y=87735 $D=8
M165 VDD 158 160 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=67235 $Y=154595 $D=8
M166 VDD 394 393 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=67235 $Y=155875 $D=8
M167 VDD 402 401 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=67235 $Y=190595 $D=8
M168 VDD 419 420 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=67235 $Y=191875 $D=8
M169 158 160 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=68375 $Y=154595 $D=8
M170 394 393 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=68375 $Y=155875 $D=8
M171 402 401 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=68375 $Y=190595 $D=8
M172 419 420 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=68375 $Y=191875 $D=8
M173 451 ypass[2] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=68145 $Y=87735 $D=8
M174 VDD 170 172 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=70235 $Y=154595 $D=8
M175 VDD 396 395 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=70235 $Y=155875 $D=8
M176 VDD 404 403 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=70235 $Y=190595 $D=8
M177 VDD 417 418 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=70235 $Y=191875 $D=8
M178 170 172 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=71375 $Y=154595 $D=8
M179 396 395 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=71375 $Y=155875 $D=8
M180 404 403 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=71375 $Y=190595 $D=8
M181 417 418 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=71375 $Y=191875 $D=8
M182 452 ypass[1] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=71810 $Y=87735 $D=8
M183 VDD 166 168 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=73235 $Y=154595 $D=8
M184 VDD 398 397 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=73235 $Y=155875 $D=8
M185 VDD 406 405 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=73235 $Y=190595 $D=8
M186 VDD 415 416 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=73235 $Y=191875 $D=8
M187 166 168 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=74375 $Y=154595 $D=8
M188 398 397 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=74375 $Y=155875 $D=8
M189 406 405 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=74375 $Y=190595 $D=8
M190 415 416 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=74375 $Y=191875 $D=8
M191 328 ypass[0] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=74340 $Y=87735 $D=8
M192 VDD 491 492 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=79235 $Y=190595 $D=8
M193 VDD 429 430 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=79235 $Y=191875 $D=8
M194 326 ypass[7] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=78015 $Y=87735 $D=8
M195 491 492 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=80375 $Y=190595 $D=8
M196 429 430 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=80375 $Y=191875 $D=8
M197 342 ypass[6] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=80540 $Y=87735 $D=8
M198 VDD 489 490 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=82235 $Y=190595 $D=8
M199 VDD 427 428 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=82235 $Y=191875 $D=8
M200 489 490 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=83375 $Y=190595 $D=8
M201 427 428 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=83375 $Y=191875 $D=8
M202 VDD 487 488 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=85235 $Y=190595 $D=8
M203 VDD 425 426 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=85235 $Y=191875 $D=8
M204 341 ypass[5] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=84205 $Y=87735 $D=8
M205 487 488 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=86375 $Y=190595 $D=8
M206 425 426 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=86375 $Y=191875 $D=8
M207 340 ypass[4] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=86735 $Y=87735 $D=8
M208 VDD 485 486 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=88235 $Y=190595 $D=8
M209 VDD 423 424 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=88235 $Y=191875 $D=8
M210 485 486 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=89375 $Y=190595 $D=8
M211 423 424 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=89375 $Y=191875 $D=8
M212 VDD 499 500 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=91235 $Y=190595 $D=8
M213 VDD 437 438 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=91235 $Y=191875 $D=8
M214 339 ypass[3] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=90395 $Y=87735 $D=8
M215 499 500 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=92375 $Y=190595 $D=8
M216 437 438 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=92375 $Y=191875 $D=8
M217 338 ypass[2] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=92925 $Y=87735 $D=8
M218 VDD 497 498 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=94235 $Y=190595 $D=8
M219 VDD 435 436 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=94235 $Y=191875 $D=8
M220 497 498 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=95375 $Y=190595 $D=8
M221 435 436 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=95375 $Y=191875 $D=8
M222 VDD 495 496 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=97235 $Y=190595 $D=8
M223 VDD 433 434 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=97235 $Y=191875 $D=8
M224 337 ypass[1] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=96590 $Y=87735 $D=8
M225 495 496 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=98375 $Y=190595 $D=8
M226 433 434 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=98375 $Y=191875 $D=8
M227 VDD 493 494 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=100235 $Y=190595 $D=8
M228 VDD 431 432 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=100235 $Y=191875 $D=8
M229 336 ypass[0] VDD VDD pmos_5p0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=99120 $Y=87735 $D=8
M230 493 494 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=101375 $Y=190595 $D=8
M231 431 432 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=101375 $Y=191875 $D=8
M232 VDD 137 138 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=106235 $Y=154595 $D=8
M233 VDD 453 454 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=106235 $Y=155875 $D=8
M234 VDD 455 456 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=106235 $Y=163595 $D=8
M235 VDD 457 458 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=106235 $Y=164875 $D=8
M236 VDD 459 460 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=106235 $Y=172595 $D=8
M237 VDD 461 462 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=106235 $Y=173875 $D=8
M238 VDD 463 464 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=106235 $Y=181595 $D=8
M239 VDD 465 466 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=106235 $Y=182875 $D=8
M240 VDD 467 468 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=106235 $Y=190595 $D=8
M241 VDD 139 140 VDD pmos_5p0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=106235 $Y=191875 $D=8
M242 VDD VSS VDD VDD pmos_5p0 L=2.365e-06 W=8.19e-05 AD=0 AS=6.1309e-11 PD=0 PS=0.000217698 NRD=0 NRS=11.8457 m=1 nf=36 $X=-3770 $Y=145970 $D=8
M243 137 138 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=107375 $Y=154595 $D=8
M244 453 454 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=107375 $Y=155875 $D=8
M245 455 456 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=107375 $Y=163595 $D=8
M246 457 458 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=107375 $Y=164875 $D=8
M247 459 460 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=107375 $Y=172595 $D=8
M248 461 462 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=107375 $Y=173875 $D=8
M249 463 464 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=107375 $Y=181595 $D=8
M250 465 466 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=107375 $Y=182875 $D=8
M251 467 468 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=107375 $Y=190595 $D=8
M252 139 140 VDD VDD pmos_5p0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=107375 $Y=191875 $D=8
X255 VSS VSS 141 142 143 144 145 146 147 148 ICV_7 $T=12605 151035 1 180 $X=9265 $Y=150695
X256 VSS VSS 149 150 151 152 153 154 155 156 ICV_7 $T=18605 151035 1 180 $X=15265 $Y=150695
X257 VSS VSS 157 158 159 160 161 162 163 164 ICV_7 $T=66605 151035 1 180 $X=63265 $Y=150695
X258 VSS VSS 165 166 167 168 169 170 171 172 ICV_7 $T=72605 151035 1 180 $X=69265 $Y=150695
X259 VSS VSS 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187 188 ICV_8 $T=605 151035 1 180 $X=-2735 $Y=150695
X260 VSS VSS 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 ICV_8 $T=605 196035 0 180 $X=-2735 $Y=191195
X261 VSS VSS 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 ICV_8 $T=12605 196035 0 180 $X=9265 $Y=191195
X262 VSS VSS 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 ICV_8 $T=27605 196035 0 180 $X=24265 $Y=191195
X263 VSS VSS 237 238 239 240 241 242 243 244 245 246 247 248 249 250 251 252 ICV_8 $T=39605 196035 0 180 $X=36265 $Y=191195
X264 VSS VSS 253 254 255 256 257 258 259 260 261 262 263 264 265 266 267 268 ICV_8 $T=54605 151035 1 180 $X=51265 $Y=150695
X275 107 VSS q[1] pcb[2] din[1] men VDD b[23] bb[23] WEN[2] b[16] bb[16] bb[17] b[17] b[18] bb[18] bb[19] b[19] b[20] bb[20]
+ bb[21] b[21] b[22] bb[22] 325 ypass[0] ypass[1] ypass[2] GWE ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] GWEN 329 330 331 332 333
+ 334 335
+ saout_R_m2 $T=51040 30 1 180 $X=12875 $Y=-18280
X276 106 VSS q[3] pcb[0] din[3] men VDD b[7] bb[7] WEN[0] b[0] bb[0] bb[1] b[1] b[2] bb[2] bb[3] b[3] b[4] bb[4]
+ bb[5] b[5] b[6] bb[6] 326 ypass[0] ypass[1] ypass[2] GWE ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] GWEN 336 337 338 339 340
+ 341 342
+ saout_R_m2 $T=105040 30 1 180 $X=66875 $Y=-18280
X277 VDD VSS WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] b[31] bb[31] bb[30] b[30] b[29] bb[29] bb[28] b[28] 343 344
+ 345 346 347 348 349 350 351 352 353 354 355 356 357 358
+ ICV_17 $T=-2395 155535 0 0 $X=-2735 $Y=155195
X278 VDD VSS WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] b[27] bb[27] bb[26] b[26] b[25] bb[25] bb[24] b[24] 359 360
+ 361 362 363 364 365 366 367 368 369 370 371 372 373 374
+ ICV_17 $T=9605 155535 0 0 $X=9265 $Y=155195
X279 VDD VSS WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] b[15] bb[15] bb[14] b[14] b[13] bb[13] bb[12] b[12] 375 376
+ 377 378 379 380 381 382 383 384 385 386 387 388 389 390
+ ICV_17 $T=51605 155535 0 0 $X=51265 $Y=155195
X280 VDD VSS WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] b[11] bb[11] bb[10] b[10] b[9] bb[9] bb[8] b[8] 391 392
+ 393 394 395 396 397 398 399 400 401 402 403 404 405 406
+ ICV_17 $T=63605 155535 0 0 $X=63265 $Y=155195
X281 VSS VSS 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422 423 424
+ 425 426 427 428 429 430 431 432 433 434 435 436 437 438
+ new_dummyrow_unit $T=51295 196920 1 0 $X=51265 $Y=191195
X282 108 VSS q[0] din[0] pcb[3] men VDD b[24] bb[24] WEN[3] b[31] bb[31] bb[30] b[30] b[29] bb[29] bb[28] b[28] b[27] bb[27]
+ bb[26] b[26] b[25] bb[25] 327 ypass[7] ypass[6] ypass[5] GWE ypass[4] ypass[3] ypass[2] ypass[1] ypass[0] GWEN 439 440 441 442 443
+ 444 445
+ saout_m2 $T=-4830 -5 0 0 $X=-6175 $Y=-17780
X283 105 VSS q[2] din[2] pcb[1] men VDD b[8] bb[8] WEN[1] b[15] bb[15] bb[14] b[14] b[13] bb[13] bb[12] b[12] b[11] bb[11]
+ bb[10] b[10] b[9] bb[9] 328 ypass[7] ypass[6] ypass[5] GWE ypass[4] ypass[3] ypass[2] ypass[1] ypass[0] GWEN 446 447 448 449 450
+ 451 452
+ saout_m2 $T=49170 -5 0 0 $X=47825 $Y=-17780
X284 46 47 VSS 453 454 455 456 ICV_25 $T=102605 160035 0 0 $X=102265 $Y=155195
X285 46 47 VSS 457 458 459 460 ICV_25 $T=102605 169035 0 0 $X=102265 $Y=164195
X286 46 47 VSS 461 462 463 464 ICV_25 $T=102605 178035 0 0 $X=102265 $Y=173195
X287 46 47 VSS 465 466 467 468 ICV_25 $T=102605 187035 0 0 $X=102265 $Y=182195
X288 VDD VSS WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] b[20] bb[20] bb[21] b[21] b[22] bb[22] bb[23] b[23] 469 470
+ 471 472 473 474 475 476
+ ICV_26 $T=27605 151035 1 180 $X=24265 $Y=150695
X289 VDD VSS WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] b[16] bb[16] bb[17] b[17] b[18] bb[18] bb[19] b[19] 477 478
+ 479 480 481 482 483 484
+ ICV_26 $T=39605 151035 1 180 $X=36265 $Y=150695
X290 VDD VSS WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] b[4] bb[4] bb[5] b[5] b[6] bb[6] bb[7] b[7] 485 486
+ 487 488 489 490 491 492
+ ICV_26 $T=81605 151035 1 180 $X=78265 $Y=150695
X291 VDD VSS WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] WL[7] b[0] bb[0] bb[1] b[1] b[2] bb[2] bb[3] b[3] 493 494
+ 495 496 497 498 499 500
+ ICV_26 $T=93605 151035 1 180 $X=90265 $Y=150695
.ENDS
***************************************
.SUBCKT M1_PSUB_CDNS_40254123696108
** N=2765 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT gf180mcu_fd_sram__64x8m8wm1 A[5] A[4] A[3] A[2] A[1] A[0] CEN CLK 
+ D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] GWEN Q[7] Q[6] Q[5] Q[4] Q[3] Q[2] 
+ Q[1] Q[0] VDD VSS WEN[7] WEN[6] WEN[5] WEN[4] WEN[3] WEN[2] WEN[1] WEN[0]
** N=5630 EP=35 IP=395 FDC=6349
M0 VSS 395 599 VSS nmos_5p0 L=6e-07 W=1.36e-06 AD=3.536e-13 AS=5.984e-13 PD=1.88e-06 PS=3.6e-06 NRD=0.191176 NRS=0.323529 m=1 nf=1 $X=233770 $Y=54135 $D=2
M1 599 CLK VSS VSS nmos_5p0 L=6e-07 W=1.36e-06 AD=5.984e-13 AS=3.536e-13 PD=3.6e-06 PS=1.88e-06 NRD=0.323529 NRS=0.191176 m=1 nf=1 $X=234890 $Y=54135 $D=2
M2 592 595 VSS VSS nmos_5p0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.58e-06 PS=1.084e-05 NRD=0.229075 NRS=0.387665 m=1 nf=2 $X=242235 $Y=54135 $D=2
M3 273 598 VSS VSS nmos_5p0 L=1e-06 W=6e-07 AD=2.64e-13 AS=2.64e-13 PD=2.08e-06 PS=2.08e-06 NRD=0.733333 NRS=0.733333 m=1 nf=1 $X=243265 $Y=46010 $D=2
M4 CEN 599 595 VSS nmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=245925 $Y=54135 $D=2
M5 242 461 VSS VSS nmos_5p0 L=6e-07 W=4.99e-05 AD=1.47704e-11 AS=1.47704e-11 PD=6.284e-05 PS=6.284e-05 NRD=0.148297 NRS=0.148297 m=1 nf=5 $X=241995 $Y=72320 $D=2
M6 309 273 VSS VSS nmos_5p0 L=6e-07 W=7.5e-07 AD=3.3e-13 AS=3.3e-13 PD=2.38e-06 PS=2.38e-06 NRD=0.586667 NRS=0.586667 m=1 nf=1 $X=246495 $Y=46075 $D=2
M7 346 309 VSS VSS nmos_5p0 L=6e-07 W=3.02e-06 AD=1.3288e-12 AS=1.3288e-12 PD=6.92e-06 PS=6.92e-06 NRD=0.145695 NRS=0.145695 m=1 nf=1 $X=249065 $Y=46070 $D=2
M8 5512 346 VSS VSS nmos_5p0 L=6e-07 W=2.268e-05 AD=5.8968e-12 AS=1.34946e-11 PD=2.32e-05 PS=4.655e-05 NRD=0.0114638 NRS=0.0262346 m=1 nf=1 $X=256125 $Y=28435 $D=2
M9 5513 CLK 5512 VSS nmos_5p0 L=6e-07 W=2.268e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=257245 $Y=28435 $D=2
M10 438 592 5513 VSS nmos_5p0 L=6e-07 W=2.268e-05 AD=1.33812e-11 AS=5.8968e-12 PD=4.654e-05 PS=2.32e-05 NRD=0.0260141 NRS=0.0114638 m=1 nf=1 $X=258365 $Y=28435 $D=2
M11 5514 488 VSS VSS nmos_5p0 L=6e-07 W=1.8145e-05 AD=4.7177e-12 AS=1.07963e-11 PD=1.8665e-05 PS=3.748e-05 NRD=0.014329 NRS=0.0327914 m=1 nf=1 $X=262120 $Y=29545 $D=2
M12 461 438 5514 VSS nmos_5p0 L=6e-07 W=1.8145e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=263240 $Y=29545 $D=2
M13 5515 438 461 VSS nmos_5p0 L=6e-07 W=1.8145e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=264360 $Y=29545 $D=2
M14 VSS 488 5515 VSS nmos_5p0 L=6e-07 W=1.8145e-05 AD=1.07055e-11 AS=4.7177e-12 PD=3.747e-05 PS=1.8665e-05 NRD=0.0325158 NRS=0.014329 m=1 nf=1 $X=265480 $Y=29545 $D=2
M15 5516 461 VSS VSS nmos_5p0 L=6e-07 W=4.54e-06 AD=1.16905e-12 AS=2.7013e-12 PD=5.055e-06 PS=1.027e-05 NRD=0.0567181 NRS=0.131057 m=1 nf=1 $X=268545 $Y=43150 $D=2
M16 488 608 5516 VSS nmos_5p0 L=6e-07 W=4.54e-06 AD=2.27e-14 AS=-2.27e-14 PD=1e-08 PS=-1e-08 NRD=0.00110132 NRS=-0.00110132 m=1 nf=1 $X=269660 $Y=43150 $D=2
M17 5517 608 488 VSS nmos_5p0 L=6e-07 W=4.54e-06 AD=-2.27e-14 AS=2.27e-14 PD=-1e-08 PS=1e-08 NRD=-0.00110132 NRS=0.00110132 m=1 nf=1 $X=270785 $Y=43150 $D=2
M18 VSS 461 5517 VSS nmos_5p0 L=6e-07 W=4.54e-06 AD=2.7013e-12 AS=1.16905e-12 PD=1.027e-05 PS=5.055e-06 NRD=0.131057 NRS=0.0567181 m=1 nf=1 $X=271900 $Y=43150 $D=2
M19 395 242 VSS VSS nmos_5p0 L=6e-07 W=0.0001474 AD=3.8324e-11 AS=4.09772e-11 PD=0.0001578 PS=0.00017326 NRD=0.705563 NRS=0.75441 m=1 nf=20 $X=253180 $Y=76320 $D=2
M20 5594 5431 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=13620 $Y=160970 $D=8
M21 5593 5431 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=13620 $Y=164845 $D=8
M22 5591 5431 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=16720 $Y=160970 $D=8
M23 5592 5431 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=16720 $Y=164845 $D=8
M24 5590 5431 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=19815 $Y=160970 $D=8
M25 5589 5431 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=19815 $Y=164845 $D=8
M26 5587 5431 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=22915 $Y=160970 $D=8
M27 5588 5431 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=22915 $Y=164845 $D=8
M28 5578 5431 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=26005 $Y=160970 $D=8
M29 5577 5431 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=26005 $Y=164845 $D=8
M30 5575 5431 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=29105 $Y=160970 $D=8
M31 5576 5431 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=29105 $Y=164845 $D=8
M32 5580 5431 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=32200 $Y=160970 $D=8
M33 5579 5431 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=32200 $Y=164845 $D=8
M34 625 5431 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=35120 $Y=160970 $D=8
M35 626 5431 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=35120 $Y=164845 $D=8
M36 627 5432 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=38575 $Y=160970 $D=8
M37 628 5432 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=38575 $Y=164845 $D=8
M38 5599 5432 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=41500 $Y=160970 $D=8
M39 5600 5432 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=41500 $Y=164845 $D=8
M40 5598 5432 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=44595 $Y=160970 $D=8
M41 5597 5432 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=44595 $Y=164845 $D=8
M42 5595 5432 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=47695 $Y=160970 $D=8
M43 5596 5432 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=47695 $Y=164845 $D=8
M44 5608 5432 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=50785 $Y=160970 $D=8
M45 5607 5432 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=50785 $Y=164845 $D=8
M46 5605 5432 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=53885 $Y=160970 $D=8
M47 5606 5432 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=53885 $Y=164845 $D=8
M48 5604 5432 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=56980 $Y=160970 $D=8
M49 5603 5432 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=56980 $Y=164845 $D=8
M50 5601 5432 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=60080 $Y=160970 $D=8
M51 5602 5432 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=60080 $Y=164845 $D=8
M52 5616 5433 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=67620 $Y=160970 $D=8
M53 5615 5433 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=67620 $Y=164845 $D=8
M54 5613 5433 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=70720 $Y=160970 $D=8
M55 5614 5433 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=70720 $Y=164845 $D=8
M56 5612 5433 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=73815 $Y=160970 $D=8
M57 5611 5433 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=73815 $Y=164845 $D=8
M58 5609 5433 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=76915 $Y=160970 $D=8
M59 5610 5433 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=76915 $Y=164845 $D=8
M60 5584 5433 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=80005 $Y=160970 $D=8
M61 5583 5433 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=80005 $Y=164845 $D=8
M62 5581 5433 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=83105 $Y=160970 $D=8
M63 5582 5433 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=83105 $Y=164845 $D=8
M64 5586 5433 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=86200 $Y=160970 $D=8
M65 5585 5433 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=86200 $Y=164845 $D=8
M66 629 5433 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=89120 $Y=160970 $D=8
M67 630 5433 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=89120 $Y=164845 $D=8
M68 631 5434 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=92575 $Y=160970 $D=8
M69 632 5434 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=92575 $Y=164845 $D=8
M70 5629 5434 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=95500 $Y=160970 $D=8
M71 5630 5434 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=95500 $Y=164845 $D=8
M72 5628 5434 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=98595 $Y=160970 $D=8
M73 5627 5434 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=98595 $Y=164845 $D=8
M74 5625 5434 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=101695 $Y=160970 $D=8
M75 5626 5434 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=101695 $Y=164845 $D=8
M76 5624 5434 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=104785 $Y=160970 $D=8
M77 5623 5434 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=104785 $Y=164845 $D=8
M78 5621 5434 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=107885 $Y=160970 $D=8
M79 5622 5434 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=107885 $Y=164845 $D=8
M80 5620 5434 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=110980 $Y=160970 $D=8
M81 5619 5434 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=110980 $Y=164845 $D=8
M82 5617 5434 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=114080 $Y=160970 $D=8
M83 5618 5434 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=114080 $Y=164845 $D=8
M84 5518 395 VDD VDD pmos_5p0 L=5.95e-07 W=2.28e-06 AD=5.985e-13 AS=1.3566e-12 PD=2.805e-06 PS=5.75e-06 NRD=0.115132 NRS=0.260965 m=1 nf=1 $X=233770 $Y=57780 $D=8
M85 593 599 VDD VDD pmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=233770 $Y=63100 $D=8
M86 599 CLK 5518 VDD pmos_5p0 L=5.95e-07 W=2.28e-06 AD=1.3566e-12 AS=5.985e-13 PD=5.75e-06 PS=2.805e-06 NRD=0.260965 NRS=0.115132 m=1 nf=1 $X=234890 $Y=57780 $D=8
M87 592 595 VDD VDD pmos_5p0 L=6e-07 W=1.134e-05 AD=2.9484e-12 AS=4.9896e-12 PD=1.238e-05 PS=2.444e-05 NRD=0.0917108 NRS=0.155203 m=1 nf=2 $X=242235 $Y=57810 $D=8
M88 273 598 VDD VDD pmos_5p0 L=1e-06 W=9e-07 AD=3.96e-13 AS=3.96e-13 PD=2.68e-06 PS=2.68e-06 NRD=0.488889 NRS=0.488889 m=1 nf=1 $X=243265 $Y=42525 $D=8
M89 CEN 593 595 VDD pmos_5p0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=245925 $Y=59010 $D=8
M90 594 599 595 VDD pmos_5p0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=245925 $Y=64875 $D=8
M91 309 273 VDD VDD pmos_5p0 L=6e-07 W=1.89e-06 AD=8.316e-13 AS=8.316e-13 PD=4.66e-06 PS=4.66e-06 NRD=0.232804 NRS=0.232804 m=1 nf=1 $X=246495 $Y=41535 $D=8
M92 346 309 VDD VDD pmos_5p0 L=6e-07 W=7.54e-06 AD=1.9604e-12 AS=3.3176e-12 PD=8.58e-06 PS=1.684e-05 NRD=0.137931 NRS=0.233422 m=1 nf=2 $X=249065 $Y=39655 $D=8
M93 242 461 VDD VDD pmos_5p0 L=6e-07 W=0.0001248 AD=3.2448e-11 AS=3.69283e-11 PD=0.00013 PS=0.000130718 NRD=0.208333 NRS=0.237099 m=1 nf=10 $X=240535 $Y=94430 $D=8
M94 438 346 VDD VDD pmos_5p0 L=6e-07 W=1.95e-05 AD=5.07e-12 AS=8.58e-12 PD=2.002e-05 PS=3.988e-05 NRD=0.0133333 NRS=0.0225641 m=1 nf=1 $X=256125 $Y=53590 $D=8
M95 VDD CLK 438 VDD pmos_5p0 L=6e-07 W=1.95e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=257245 $Y=53590 $D=8
M96 438 592 VDD VDD pmos_5p0 L=6e-07 W=1.95e-05 AD=8.58e-12 AS=5.07e-12 PD=3.988e-05 PS=2.002e-05 NRD=0.0225641 NRS=0.0133333 m=1 nf=1 $X=258365 $Y=53590 $D=8
M97 VDD 488 461 VDD pmos_5p0 L=6e-07 W=2.268e-05 AD=5.8968e-12 AS=9.9792e-12 PD=2.32e-05 PS=4.624e-05 NRD=0.0114638 NRS=0.0194004 m=1 nf=1 $X=262120 $Y=50420 $D=8
M98 461 438 VDD VDD pmos_5p0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.64e-05 PS=4.64e-05 NRD=0.0229277 NRS=0.0229277 m=1 nf=2 $X=263240 $Y=50420 $D=8
M99 461 488 VDD VDD pmos_5p0 L=6e-07 W=2.268e-05 AD=9.9792e-12 AS=5.8968e-12 PD=4.624e-05 PS=2.32e-05 NRD=0.0194004 NRS=0.0114638 m=1 nf=1 $X=265480 $Y=50420 $D=8
M100 VDD 461 488 VDD pmos_5p0 L=6e-07 W=2.268e-05 AD=5.8968e-12 AS=9.9792e-12 PD=2.32e-05 PS=4.624e-05 NRD=0.0114638 NRS=0.0194004 m=1 nf=1 $X=268545 $Y=50420 $D=8
M101 488 608 VDD VDD pmos_5p0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.64e-05 PS=4.64e-05 NRD=0.0229277 NRS=0.0229277 m=1 nf=2 $X=269665 $Y=50420 $D=8
M102 488 461 VDD VDD pmos_5p0 L=6e-07 W=2.268e-05 AD=9.9792e-12 AS=5.8968e-12 PD=4.624e-05 PS=2.32e-05 NRD=0.0194004 NRS=0.0114638 m=1 nf=1 $X=271905 $Y=50420 $D=8
M103 395 242 VDD VDD pmos_5p0 L=6e-07 W=0.0003674 AD=9.5524e-11 AS=1.02119e-10 PD=0.0003778 PS=0.000378518 NRD=0.28307 NRS=0.302613 m=1 nf=20 $X=253180 $Y=88540 $D=8
M104 5566 5428 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=311500 $Y=160970 $D=8
M105 5565 5428 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=311500 $Y=164845 $D=8
M106 5563 5428 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=314600 $Y=160970 $D=8
M107 5564 5428 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=314600 $Y=164845 $D=8
M108 5562 5428 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=317695 $Y=160970 $D=8
M109 5561 5428 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=317695 $Y=164845 $D=8
M110 5559 5428 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=320795 $Y=160970 $D=8
M111 5560 5428 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=320795 $Y=164845 $D=8
M112 5550 5428 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=323885 $Y=160970 $D=8
M113 5549 5428 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=323885 $Y=164845 $D=8
M114 5547 5428 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=326985 $Y=160970 $D=8
M115 5548 5428 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=326985 $Y=164845 $D=8
M116 5552 5428 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=330080 $Y=160970 $D=8
M117 5551 5428 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=330080 $Y=164845 $D=8
M118 617 5428 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=333000 $Y=160970 $D=8
M119 618 5428 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=333000 $Y=164845 $D=8
M120 619 5429 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=336455 $Y=160970 $D=8
M121 620 5429 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=336455 $Y=164845 $D=8
M122 5523 5429 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=339380 $Y=160970 $D=8
M123 5524 5429 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=339380 $Y=164845 $D=8
M124 5522 5429 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=342475 $Y=160970 $D=8
M125 5521 5429 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=342475 $Y=164845 $D=8
M126 5519 5429 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=345575 $Y=160970 $D=8
M127 5520 5429 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=345575 $Y=164845 $D=8
M128 5532 5429 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=348665 $Y=160970 $D=8
M129 5531 5429 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=348665 $Y=164845 $D=8
M130 5529 5429 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=351765 $Y=160970 $D=8
M131 5530 5429 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=351765 $Y=164845 $D=8
M132 5528 5429 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=354860 $Y=160970 $D=8
M133 5527 5429 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=354860 $Y=164845 $D=8
M134 5525 5429 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=357960 $Y=160970 $D=8
M135 5526 5429 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=357960 $Y=164845 $D=8
M136 5574 5430 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=365500 $Y=160970 $D=8
M137 5573 5430 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=365500 $Y=164845 $D=8
M138 5571 5430 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=368600 $Y=160970 $D=8
M139 5572 5430 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=368600 $Y=164845 $D=8
M140 5570 5430 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=371695 $Y=160970 $D=8
M141 5569 5430 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=371695 $Y=164845 $D=8
M142 5567 5430 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=374795 $Y=160970 $D=8
M143 5568 5430 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=374795 $Y=164845 $D=8
M144 5556 5430 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=377885 $Y=160970 $D=8
M145 5555 5430 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=377885 $Y=164845 $D=8
M146 5553 5430 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=380985 $Y=160970 $D=8
M147 5554 5430 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=380985 $Y=164845 $D=8
M148 5558 5430 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=384080 $Y=160970 $D=8
M149 5557 5430 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=384080 $Y=164845 $D=8
M150 621 5430 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=387000 $Y=160970 $D=8
M151 622 5430 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=387000 $Y=164845 $D=8
M152 623 616 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=390455 $Y=160970 $D=8
M153 624 616 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=390455 $Y=164845 $D=8
M154 5537 616 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=393380 $Y=160970 $D=8
M155 5538 616 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=393380 $Y=164845 $D=8
M156 5536 616 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=396475 $Y=160970 $D=8
M157 5535 616 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=396475 $Y=164845 $D=8
M158 5533 616 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=399575 $Y=160970 $D=8
M159 5534 616 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=399575 $Y=164845 $D=8
M160 5546 616 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=402665 $Y=160970 $D=8
M161 5545 616 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=402665 $Y=164845 $D=8
M162 5543 616 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=405765 $Y=160970 $D=8
M163 5544 616 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=405765 $Y=164845 $D=8
M164 5542 616 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=408860 $Y=160970 $D=8
M165 5541 616 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=408860 $Y=164845 $D=8
M166 5539 616 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=411960 $Y=160970 $D=8
M167 5540 616 VDD VDD pmos_5p0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=411960 $Y=164845 $D=8
X175 VSS 593 599 VSS nmos_1p2$$46563372 $T=233925 66830 0 0 $X=232780 $Y=66145
X176 594 VSS 592 VSS nmos_1p2$$46563372 $T=243510 68190 1 0 $X=242365 $Y=66555
X177 595 594 593 VSS nmos_1p2$$46563372 $T=246080 68190 1 0 $X=244935 $Y=66555
X178 VDD 594 592 pmos_1p2$$46273580 $T=242390 65835 1 0 $X=240960 $Y=64015
X180 VSS 608 616 VDD 5452 WEN[5] 5429 619 620 395 WEN[7] 623 624 WEN[4] 5428 617 618 WEN[6] 5430 621
+ 622 5461 5462 5463 5464 5465 5466 5467 5468 607 5451 5459 5460 5458 5457 5456 5455 5454 5453 D[5]
+ Q[5] D[7] Q[7] D[4] Q[4] D[6] Q[6] 5519 5520 5521 5522 5523 5524 5525 5526 5527 5528 5529 5530 5531
+ 5532 5533 5534 5535 5536 5537 5538 5539 5540 5541 5542 5543 5544 5545 5546 5547 5548 5549 5550 5551
+ 5552 5553 5554 5555 5556 5557 5558 5559 5560 5561 5562 5563 5564 5565 5566 5567 5568 5569 5570 5571
+ 5572 5573 5574
+ rcol4_64 $T=302555 25095 0 0 $X=297105 $Y=5955
X191 VSS 597 CLK nmos_5p0_CDNS_4025412369694 $T=234280 46585 1 0 $X=233600 $Y=45365
X192 VSS 598 597 nmos_5p0_CDNS_4025412369694 $T=239670 46585 1 0 $X=238990 $Y=45365
X193 VDD 597 CLK pmos_5p0_CDNS_4025412369691 $T=234280 43425 1 0 $X=233240 $Y=41905
X194 VDD 598 597 pmos_5p0_CDNS_4025412369691 $T=239670 43425 1 0 $X=238630 $Y=41905
X197 VSS 395 VDD CLK A[5] A[4] A[3] 5496 5497 5498 5499 5500 5501 5502 5503 xpredec1 $T=219860 111460 0 0 $X=219855 $Y=111455
X198 VSS 5450 VDD GWEN CLK 5451 607 wen_v2 $T=208415 16605 0 0 $X=208280 $Y=15275
X201 VSS VDD 395 CLK VSS VSS 5485 5486 5490 5491 xpredec0 $T=146075 111460 0 0 $X=144630 $Y=111455
X202 VSS VDD 395 CLK VSS VSS 5492 5493 5494 5495 xpredec0 $T=182970 111460 0 0 $X=181525 $Y=111455
X203 VSS VDD 395 CLK 5448 5449 5442 5443 5444 5445 5446 5447 5460 5459 5458 5457 5456 5455 5454 5453
+ A[2] A[1] A[0]
+ ypredec1 $T=145470 26355 0 0 $X=146365 $Y=26735
X205 395 VSS 5452 VDD 5503 5502 5501 5500 5499 5498 5497 5496 5469 5470 5471 5472 5473 5474 5475 5476
+ 5462 5463 5465 5467 5468 5464 5466 5461
+ xdec8_64 $T=143385 180635 0 0 $X=126565 $Y=178920
X206 VSS VDD WEN[1] 5432 627 628 395 WEN[3] 5434 631 632 WEN[0] 5431 625 626 WEN[2] 5433 629 630 5469
+ 5470 5471 5472 5473 5474 5475 5476 5451 607 5442 5443 5444 5445 5446 5447 5448 5449 D[1] Q[1] D[3]
+ Q[3] D[0] Q[0] D[2] Q[2] 5575 5576 5577 5578 5579 5580 5581 5582 5583 5584 5585 5586 5587 5588 5589
+ 5590 5591 5592 5593 5594 5595 5596 5597 5598 5599 5600 5601 5602 5603 5604 5605 5606 5607 5608 5609
+ 5610 5611 5612 5613 5614 5615 5616 5617 5618 5619 5620 5621 5622 5623 5624 5625 5626 5627 5628 5629
+ 5630
+ lcol4_64 $T=14605 25095 0 0 $X=2855 $Y=4030
.ENDS
***************************************
