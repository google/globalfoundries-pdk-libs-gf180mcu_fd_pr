*Xyce Common Source Circuit
** library calling


*****************
** main netlist
*****************
Vn n 0 DC 1

xrn n 0 {{device}} L={{width}}u W={{length}}u


*****************
** Analysis
*****************
.OP
.STEP TEMP {{temp}} -60 200
.print DC FORMAT=CSV file={{device}}_r_{{corner}}_temp/simulated_r/{{i}}_simulated_w{{width}}_l{{length}}.csv {(V(n)*{{length}}u)/(-I(Vn)*{{width}}u)}



.include "../../../../../design.xyce"
.lib "../../../../../sm141064.xyce" res_{{corner}}

.end