*****
***** Welcome to the Xyce(TM) Parallel Electronic Simulator
*****
***** This is version Xyce Release 7.6-opensource


** library calling

.include "../../../design.xyce"
.lib "../../../sm141064.xyce" typical

vds D_tn 0 dc 0
vgs G_tn 0 dc 3.3
vbs S_tn 0 dc 0


* circuit
xmn1 D_tn G_tn 0 S_tn {{device}} W = {{width}}u L = {{length}}u nf={{nf}} ad={{AD}}u pd={{PD}}u as={{AS}}u ps={{PS}}u TEMP=25



* measurement setup 
.meas tran vds1 AVG v(D_tn) FROM=0.1ns TO=0.2ns

* simulation setup
.tran 1ns 4ns 0.5ns

* print setup
.print tran vds1
.end