***************************
** nfet_10v0_asym_id
***************************
* Copyright 2023 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

vds D_tn 0 dc {{vds_val}}
vgs G_tn 0 dc 10
Vbs B_tn 0 dc {{vbs_val}}

.STEP TEMP {{temp}} {{temp}} {{temp}}

xmn1 D_tn G_tn 0 B_tn {{device}} W = {{width}}u L = {{length}}u

**** begin architecture code
.DC {{sweeps}}

.print DC FORMAT=CSV file={{result_path}} v(D_tn) v(G_tn) v(B_tn) {-I(Vds)}

** library calling

.include {{model_design_path}}
.lib {{model_card_path}} {{corner}}

**** end architecture code

.end
