************************************************************************
* auCdl Netlist:
* 
* Library Name:  TCG_Library
* Top Cell Name: cap_mim_1f0_m2m3_noshield
* View Name:     schematic
* Netlisted on:  Nov 24 10:39:22 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: TCG_Library
* Cell Name:    cap_mim_1f0_m2m3_noshield
* View Name:    schematic
************************************************************************

.SUBCKT cap_mim_1f0_m2m3_noshield I1_0_0_R0_BOT I1_0_0_R0_TOP I1_0_1_R0_BOT I1_0_1_R0_TOP 
+ I1_0_2_R0_BOT I1_0_2_R0_TOP I1_1_0_R0_BOT I1_1_0_R0_TOP I1_1_1_R0_BOT 
+ I1_1_1_R0_TOP I1_1_2_R0_BOT I1_1_2_R0_TOP I1_2_0_R0_BOT I1_2_0_R0_TOP 
+ I1_2_1_R0_BOT I1_2_1_R0_TOP I1_2_2_R0_BOT I1_2_2_R0_TOP I1_default_BOT 
+ I1_default_TOP
*.PININFO I1_0_0_R0_BOT:I I1_0_0_R0_TOP:I I1_0_1_R0_BOT:I I1_0_1_R0_TOP:I 
*.PININFO I1_0_2_R0_BOT:I I1_0_2_R0_TOP:I I1_1_0_R0_BOT:I I1_1_0_R0_TOP:I 
*.PININFO I1_1_1_R0_BOT:I I1_1_1_R0_TOP:I I1_1_2_R0_BOT:I I1_1_2_R0_TOP:I 
*.PININFO I1_2_0_R0_BOT:I I1_2_0_R0_TOP:I I1_2_1_R0_BOT:I I1_2_1_R0_TOP:I 
*.PININFO I1_2_2_R0_BOT:I I1_2_2_R0_TOP:I I1_default_BOT:I I1_default_TOP:I
CI1_2_2_R0 I1_2_2_R0_TOP I1_2_2_R0_BOT $[cap_mim_1f0_m2m3_noshield] M=1 l=50.000u w=50.000u 
+ c=2.5335p
CI1_2_1_R0 I1_2_1_R0_TOP I1_2_1_R0_BOT $[cap_mim_1f0_m2m3_noshield] M=1 l=50.000u w=11.560u 
+ c=0.6111156p
CI1_2_0_R0 I1_2_0_R0_TOP I1_2_0_R0_BOT $[cap_mim_1f0_m2m3_noshield] M=1 l=50.000u w=5.000u 
+ c=0.28305p
CI1_1_2_R0 I1_1_2_R0_TOP I1_1_2_R0_BOT $[cap_mim_1f0_m2m3_noshield] M=1 l=11.560u w=50.000u 
+ c=0.6111156p
CI1_1_1_R0 I1_1_1_R0_TOP I1_1_1_R0_BOT $[cap_mim_1f0_m2m3_noshield] M=1 l=11.560u w=11.560u 
+ c=0.14715556p
CI1_1_0_R0 I1_1_0_R0_TOP I1_1_0_R0_BOT $[cap_mim_1f0_m2m3_noshield] M=1 l=11.560u w=5.000u 
+ c=0.0679782p
CI1_0_2_R0 I1_0_2_R0_TOP I1_0_2_R0_BOT $[cap_mim_1f0_m2m3_noshield] M=1 l=5.000u w=50.000u 
+ c=0.28305p
CI1_0_1_R0 I1_0_1_R0_TOP I1_0_1_R0_BOT $[cap_mim_1f0_m2m3_noshield] M=1 l=5.000u w=11.560u 
+ c=0.0679782p
CI1_0_0_R0 I1_0_0_R0_TOP I1_0_0_R0_BOT $[cap_mim_1f0_m2m3_noshield] M=1 l=5.000u w=5.000u 
+ c=0.031275p
CI1_default I1_default_TOP I1_default_BOT $[cap_mim_1f0_m2m3_noshield] M=1 l=5u w=5u 
+ c=0.031275p
.ENDS

