*****************
** main netlist
*****************

Vcp c 0 dc -3
Ib f b -9u
Vbb 0 f dc=0
.temp {{temp}}
.options tnom={{temp}}

xq1 c b 0 {{device}}


*****************
** Analysis
*****************

.control
set filetype=ascii
set wr_singlescale
set wr_vecnames
dc Vcp 0 -3 -0.1 Ib -1u -9u -2u

wrdata bjt_iv_regr/pnp/ib_simulated/simulated_{{device}}_t{{temp}}.csv i(Vcp) i(Vbb)
.endc

.include "../../../design.ngspice"
.lib "../../../sm141064.ngspice" bjt_typical



.end
