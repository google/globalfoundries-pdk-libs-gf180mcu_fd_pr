
xmn1 D_tn G_tn 0 0 {{device}} W={{width}}u L={{length}}u ad={{AD}}u pd={{PD}}u as={{AS}}u ps={{PS}}u

*****************
** Analysis
*****************
.DC Vds {{vds}} Vgs {{vgs}}
.STEP TEMP {{temp}} -60 200
.print DC FORMAT=CSV file=mos_iv_reg/{{device}}/{{device}}_netlists_Rds/t{{temp}}_simulated_W{{width}}_L{{length}}.csv {1/N(xmn1:m0:gds)} v(D_tn) v(G_tn)

.include "../../../../../../design.xyce"
.lib "../../../../../../sm141064.xyce" typical

.end


* ***************************
* ** pfet_03v3_t_Rds
* ***************************
* * Copyright 2023 Efabless Corporation
* *
* * Licensed under the Apache License, Version 2.0 (the "License");
* * you may not use this file except in compliance with the License.
* * You may obtain a copy of the License at
* *
* *      http://www.apache.org/licenses/LICENSE-2.0
* *
* * Unless required by applicable law or agreed to in writing, software
* * distributed under the License is distributed on an "AS IS" BASIS,
* * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* * See the License for the specific language governing permissions and
* * limitations under the License.

vds D_tn 0 dc {{vds_val}}
vgs G_tn 0 dc -3.3
Vbs B_tn 0 dc {{vbs_val}}

.STEP TEMP {{temp}} -60 200

xmp1 D_tn G_tn 0 B_tn {{device}} W = {{width}}u L = {{length}}u

**** begin architecture code
.DC {{sweeps}}

** Get all voltages and currrent

.print DC FORMAT=CSV file={{result_path}} v(D_tn) v(G_tn) v(B_tn) {1/N(xmp1:m0:gds)} 

** library calling

.include {{model_design_path}}
.lib {{model_card_path}} {{corner}}

**** end architecture code

.end
