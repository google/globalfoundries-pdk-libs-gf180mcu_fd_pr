************************************************************************
* auCdl Netlist:
* 
* Library Name:  TCG_Library
* Top Cell Name: diode_nd2ps_03v3_dn
* View Name:     schematic
* Netlisted on:  Nov 24 09:17:22 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: TCG_Library
* Cell Name:    diode_nd2ps_03v3_dn
* View Name:    schematic
************************************************************************

.SUBCKT diode_nd2ps_03v3_dn I1_0_0_0_0_R0_MINUS I1_0_0_0_0_R0_PLUS I1_0_1_0_0_R0_MINUS 
+ I1_0_1_0_0_R0_PLUS I1_0_2_0_0_R0_MINUS I1_0_2_0_0_R0_PLUS 
+ I1_0_3_0_0_R0_MINUS I1_0_3_0_0_R0_PLUS I1_1_0_0_0_R0_MINUS 
+ I1_1_0_0_0_R0_PLUS I1_1_1_0_0_R0_MINUS I1_1_1_0_0_R0_PLUS 
+ I1_1_2_0_0_R0_MINUS I1_1_2_0_0_R0_PLUS I1_1_3_0_0_R0_MINUS 
+ I1_1_3_0_0_R0_PLUS I1_2_0_0_0_R0_MINUS I1_2_0_0_0_R0_PLUS 
+ I1_2_1_0_0_R0_MINUS I1_2_1_0_0_R0_PLUS I1_2_2_0_0_R0_MINUS 
+ I1_2_2_0_0_R0_PLUS I1_2_3_0_0_R0_MINUS I1_2_3_0_0_R0_PLUS 
+ I1_3_0_0_0_R0_MINUS I1_3_0_0_0_R0_PLUS I1_3_1_0_0_R0_MINUS 
+ I1_3_1_0_0_R0_PLUS I1_3_2_0_0_R0_MINUS I1_3_2_0_0_R0_PLUS 
+ I1_3_3_0_0_R0_MINUS I1_3_3_0_0_R0_PLUS I1_default_MINUS I1_default_PLUS
*.PININFO I1_0_0_0_0_R0_MINUS:I I1_0_0_0_0_R0_PLUS:I I1_0_1_0_0_R0_MINUS:I 
*.PININFO I1_0_1_0_0_R0_PLUS:I I1_0_2_0_0_R0_MINUS:I I1_0_2_0_0_R0_PLUS:I 
*.PININFO I1_0_3_0_0_R0_MINUS:I I1_0_3_0_0_R0_PLUS:I I1_1_0_0_0_R0_MINUS:I 
*.PININFO I1_1_0_0_0_R0_PLUS:I I1_1_1_0_0_R0_MINUS:I I1_1_1_0_0_R0_PLUS:I 
*.PININFO I1_1_2_0_0_R0_MINUS:I I1_1_2_0_0_R0_PLUS:I I1_1_3_0_0_R0_MINUS:I 
*.PININFO I1_1_3_0_0_R0_PLUS:I I1_2_0_0_0_R0_MINUS:I I1_2_0_0_0_R0_PLUS:I 
*.PININFO I1_2_1_0_0_R0_MINUS:I I1_2_1_0_0_R0_PLUS:I I1_2_2_0_0_R0_MINUS:I 
*.PININFO I1_2_2_0_0_R0_PLUS:I I1_2_3_0_0_R0_MINUS:I I1_2_3_0_0_R0_PLUS:I 
*.PININFO I1_3_0_0_0_R0_MINUS:I I1_3_0_0_0_R0_PLUS:I I1_3_1_0_0_R0_MINUS:I 
*.PININFO I1_3_1_0_0_R0_PLUS:I I1_3_2_0_0_R0_MINUS:I I1_3_2_0_0_R0_PLUS:I 
*.PININFO I1_3_3_0_0_R0_MINUS:I I1_3_3_0_0_R0_PLUS:I I1_default_MINUS:I 
*.PININFO I1_default_PLUS:I
DI1_3_3_0_0_R0 I1_3_3_0_0_R0_PLUS I1_3_3_0_0_R0_MINUS diode_nd2ps_03v3_dn m=1 AREA=10n 
+ PJ=400u
DI1_3_2_0_0_R0 I1_3_2_0_0_R0_PLUS I1_3_2_0_0_R0_MINUS diode_nd2ps_03v3_dn m=1 AREA=1.32n 
+ PJ=226.4u
DI1_3_1_0_0_R0 I1_3_1_0_0_R0_PLUS I1_3_1_0_0_R0_MINUS diode_nd2ps_03v3_dn m=1 AREA=110p 
+ PJ=202.2u
DI1_3_0_0_0_R0 I1_3_0_0_0_R0_PLUS I1_3_0_0_0_R0_MINUS diode_nd2ps_03v3_dn m=1 AREA=56.5p 
+ PJ=201.13u
DI1_2_3_0_0_R0 I1_2_3_0_0_R0_PLUS I1_2_3_0_0_R0_MINUS diode_nd2ps_03v3_dn m=1 AREA=1.32n 
+ PJ=226.4u
DI1_2_2_0_0_R0 I1_2_2_0_0_R0_PLUS I1_2_2_0_0_R0_MINUS diode_nd2ps_03v3_dn m=1 
+ AREA=174.24p PJ=52.8u
DI1_2_1_0_0_R0 I1_2_1_0_0_R0_PLUS I1_2_1_0_0_R0_MINUS diode_nd2ps_03v3_dn m=1 
+ AREA=14.52p PJ=28.6u
DI1_2_0_0_0_R0 I1_2_0_0_0_R0_PLUS I1_2_0_0_0_R0_MINUS diode_nd2ps_03v3_dn m=1 
+ AREA=7.458p PJ=27.53u
DI1_1_3_0_0_R0 I1_1_3_0_0_R0_PLUS I1_1_3_0_0_R0_MINUS diode_nd2ps_03v3_dn m=1 AREA=110p 
+ PJ=202.2u
DI1_1_2_0_0_R0 I1_1_2_0_0_R0_PLUS I1_1_2_0_0_R0_MINUS diode_nd2ps_03v3_dn m=1 
+ AREA=14.52p PJ=28.6u
DI1_1_1_0_0_R0 I1_1_1_0_0_R0_PLUS I1_1_1_0_0_R0_MINUS diode_nd2ps_03v3_dn m=1 AREA=1.21p 
+ PJ=4.4u
DI1_1_0_0_0_R0 I1_1_0_0_0_R0_PLUS I1_1_0_0_0_R0_MINUS diode_nd2ps_03v3_dn m=1 
+ AREA=621.5f PJ=3.33u
DI1_0_3_0_0_R0 I1_0_3_0_0_R0_PLUS I1_0_3_0_0_R0_MINUS diode_nd2ps_03v3_dn m=1 AREA=56.5p 
+ PJ=201.13u
DI1_0_2_0_0_R0 I1_0_2_0_0_R0_PLUS I1_0_2_0_0_R0_MINUS diode_nd2ps_03v3_dn m=1 
+ AREA=7.458p PJ=27.53u
DI1_0_1_0_0_R0 I1_0_1_0_0_R0_PLUS I1_0_1_0_0_R0_MINUS diode_nd2ps_03v3_dn m=1 
+ AREA=621.5f PJ=3.33u
DI1_0_0_0_0_R0 I1_0_0_0_0_R0_PLUS I1_0_0_0_0_R0_MINUS diode_nd2ps_03v3_dn m=1 
+ AREA=319.225f PJ=2.26u
DI1_default I1_default_PLUS I1_default_MINUS diode_nd2ps_03v3_dn m=1 AREA=1p PJ=4u
.ENDS

