************************************************************************
* auCdl Netlist:
* 
* Library Name:  TCG_Library
* Top Cell Name: pplus_u
* View Name:     schematic
* Netlisted on:  Nov 24 09:54:02 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL gnd!

*.PIN gnd!

************************************************************************
* Library Name: TCG_Library
* Cell Name:    pplus_u
* View Name:    schematic
************************************************************************

.SUBCKT pplus_u I1_0_0_0_0_0_R0_MINUS I1_0_0_0_0_0_R0_PLUS 
+ I1_0_0_0_1_0_R0_MINUS I1_0_0_0_1_0_R0_PLUS I1_0_0_1_0_0_R0_MINUS 
+ I1_0_0_1_0_0_R0_PLUS I1_0_0_1_1_0_R0_MINUS I1_0_0_1_1_0_R0_PLUS 
+ I1_0_0_2_0_0_R0_MINUS I1_0_0_2_0_0_R0_PLUS I1_0_0_2_1_0_R0_MINUS 
+ I1_0_0_2_1_0_R0_PLUS I1_0_1_0_0_0_R0_MINUS I1_0_1_0_0_0_R0_PLUS 
+ I1_0_1_0_1_0_R0_MINUS I1_0_1_0_1_0_R0_PLUS I1_0_1_1_0_0_R0_MINUS 
+ I1_0_1_1_0_0_R0_PLUS I1_0_1_1_1_0_R0_MINUS I1_0_1_1_1_0_R0_PLUS 
+ I1_0_1_2_0_0_R0_MINUS I1_0_1_2_0_0_R0_PLUS I1_0_1_2_1_0_R0_MINUS 
+ I1_0_1_2_1_0_R0_PLUS I1_0_2_0_0_0_R0_MINUS I1_0_2_0_0_0_R0_PLUS 
+ I1_0_2_0_1_0_R0_MINUS I1_0_2_0_1_0_R0_PLUS I1_0_2_1_0_0_R0_MINUS 
+ I1_0_2_1_0_0_R0_PLUS I1_0_2_1_1_0_R0_MINUS I1_0_2_1_1_0_R0_PLUS 
+ I1_0_2_2_0_0_R0_MINUS I1_0_2_2_0_0_R0_PLUS I1_0_2_2_1_0_R0_MINUS 
+ I1_0_2_2_1_0_R0_PLUS I1_1_0_0_0_0_R0_MINUS I1_1_0_0_0_0_R0_PLUS 
+ I1_1_0_0_1_0_R0_MINUS I1_1_0_0_1_0_R0_PLUS I1_1_0_1_0_0_R0_MINUS 
+ I1_1_0_1_0_0_R0_PLUS I1_1_0_1_1_0_R0_MINUS I1_1_0_1_1_0_R0_PLUS 
+ I1_1_0_2_0_0_R0_MINUS I1_1_0_2_0_0_R0_PLUS I1_1_0_2_1_0_R0_MINUS 
+ I1_1_0_2_1_0_R0_PLUS I1_1_1_0_0_0_R0_MINUS I1_1_1_0_0_0_R0_PLUS 
+ I1_1_1_0_1_0_R0_MINUS I1_1_1_0_1_0_R0_PLUS I1_1_1_1_0_0_R0_MINUS 
+ I1_1_1_1_0_0_R0_PLUS I1_1_1_1_1_0_R0_MINUS I1_1_1_1_1_0_R0_PLUS 
+ I1_1_1_2_0_0_R0_MINUS I1_1_1_2_0_0_R0_PLUS I1_1_1_2_1_0_R0_MINUS 
+ I1_1_1_2_1_0_R0_PLUS I1_1_2_0_0_0_R0_MINUS I1_1_2_0_0_0_R0_PLUS 
+ I1_1_2_0_1_0_R0_MINUS I1_1_2_0_1_0_R0_PLUS I1_1_2_1_0_0_R0_MINUS 
+ I1_1_2_1_0_0_R0_PLUS I1_1_2_1_1_0_R0_MINUS I1_1_2_1_1_0_R0_PLUS 
+ I1_1_2_2_0_0_R0_MINUS I1_1_2_2_0_0_R0_PLUS I1_1_2_2_1_0_R0_MINUS 
+ I1_1_2_2_1_0_R0_PLUS I1_2_0_0_0_0_R0_MINUS I1_2_0_0_0_0_R0_PLUS 
+ I1_2_0_0_1_0_R0_MINUS I1_2_0_0_1_0_R0_PLUS I1_2_0_1_0_0_R0_MINUS 
+ I1_2_0_1_0_0_R0_PLUS I1_2_0_1_1_0_R0_MINUS I1_2_0_1_1_0_R0_PLUS 
+ I1_2_0_2_0_0_R0_MINUS I1_2_0_2_0_0_R0_PLUS I1_2_0_2_1_0_R0_MINUS 
+ I1_2_0_2_1_0_R0_PLUS I1_2_1_0_0_0_R0_MINUS I1_2_1_0_0_0_R0_PLUS 
+ I1_2_1_0_1_0_R0_MINUS I1_2_1_0_1_0_R0_PLUS I1_2_1_1_0_0_R0_MINUS 
+ I1_2_1_1_0_0_R0_PLUS I1_2_1_1_1_0_R0_MINUS I1_2_1_1_1_0_R0_PLUS 
+ I1_2_1_2_0_0_R0_MINUS I1_2_1_2_0_0_R0_PLUS I1_2_1_2_1_0_R0_MINUS 
+ I1_2_1_2_1_0_R0_PLUS I1_2_2_0_0_0_R0_MINUS I1_2_2_0_0_0_R0_PLUS 
+ I1_2_2_0_1_0_R0_MINUS I1_2_2_0_1_0_R0_PLUS I1_2_2_1_0_0_R0_MINUS 
+ I1_2_2_1_0_0_R0_PLUS I1_2_2_1_1_0_R0_MINUS I1_2_2_1_1_0_R0_PLUS 
+ I1_2_2_2_0_0_R0_MINUS I1_2_2_2_0_0_R0_PLUS I1_2_2_2_1_0_R0_MINUS 
+ I1_2_2_2_1_0_R0_PLUS I1_default_MINUS I1_default_PLUS gnd!
*.PININFO I1_0_0_0_0_0_R0_MINUS:I I1_0_0_0_0_0_R0_PLUS:I 
*.PININFO I1_0_0_0_1_0_R0_MINUS:I I1_0_0_0_1_0_R0_PLUS:I 
*.PININFO I1_0_0_1_0_0_R0_MINUS:I I1_0_0_1_0_0_R0_PLUS:I 
*.PININFO I1_0_0_1_1_0_R0_MINUS:I I1_0_0_1_1_0_R0_PLUS:I 
*.PININFO I1_0_0_2_0_0_R0_MINUS:I I1_0_0_2_0_0_R0_PLUS:I 
*.PININFO I1_0_0_2_1_0_R0_MINUS:I I1_0_0_2_1_0_R0_PLUS:I 
*.PININFO I1_0_1_0_0_0_R0_MINUS:I I1_0_1_0_0_0_R0_PLUS:I 
*.PININFO I1_0_1_0_1_0_R0_MINUS:I I1_0_1_0_1_0_R0_PLUS:I 
*.PININFO I1_0_1_1_0_0_R0_MINUS:I I1_0_1_1_0_0_R0_PLUS:I 
*.PININFO I1_0_1_1_1_0_R0_MINUS:I I1_0_1_1_1_0_R0_PLUS:I 
*.PININFO I1_0_1_2_0_0_R0_MINUS:I I1_0_1_2_0_0_R0_PLUS:I 
*.PININFO I1_0_1_2_1_0_R0_MINUS:I I1_0_1_2_1_0_R0_PLUS:I 
*.PININFO I1_0_2_0_0_0_R0_MINUS:I I1_0_2_0_0_0_R0_PLUS:I 
*.PININFO I1_0_2_0_1_0_R0_MINUS:I I1_0_2_0_1_0_R0_PLUS:I 
*.PININFO I1_0_2_1_0_0_R0_MINUS:I I1_0_2_1_0_0_R0_PLUS:I 
*.PININFO I1_0_2_1_1_0_R0_MINUS:I I1_0_2_1_1_0_R0_PLUS:I 
*.PININFO I1_0_2_2_0_0_R0_MINUS:I I1_0_2_2_0_0_R0_PLUS:I 
*.PININFO I1_0_2_2_1_0_R0_MINUS:I I1_0_2_2_1_0_R0_PLUS:I 
*.PININFO I1_1_0_0_0_0_R0_MINUS:I I1_1_0_0_0_0_R0_PLUS:I 
*.PININFO I1_1_0_0_1_0_R0_MINUS:I I1_1_0_0_1_0_R0_PLUS:I 
*.PININFO I1_1_0_1_0_0_R0_MINUS:I I1_1_0_1_0_0_R0_PLUS:I 
*.PININFO I1_1_0_1_1_0_R0_MINUS:I I1_1_0_1_1_0_R0_PLUS:I 
*.PININFO I1_1_0_2_0_0_R0_MINUS:I I1_1_0_2_0_0_R0_PLUS:I 
*.PININFO I1_1_0_2_1_0_R0_MINUS:I I1_1_0_2_1_0_R0_PLUS:I 
*.PININFO I1_1_1_0_0_0_R0_MINUS:I I1_1_1_0_0_0_R0_PLUS:I 
*.PININFO I1_1_1_0_1_0_R0_MINUS:I I1_1_1_0_1_0_R0_PLUS:I 
*.PININFO I1_1_1_1_0_0_R0_MINUS:I I1_1_1_1_0_0_R0_PLUS:I 
*.PININFO I1_1_1_1_1_0_R0_MINUS:I I1_1_1_1_1_0_R0_PLUS:I 
*.PININFO I1_1_1_2_0_0_R0_MINUS:I I1_1_1_2_0_0_R0_PLUS:I 
*.PININFO I1_1_1_2_1_0_R0_MINUS:I I1_1_1_2_1_0_R0_PLUS:I 
*.PININFO I1_1_2_0_0_0_R0_MINUS:I I1_1_2_0_0_0_R0_PLUS:I 
*.PININFO I1_1_2_0_1_0_R0_MINUS:I I1_1_2_0_1_0_R0_PLUS:I 
*.PININFO I1_1_2_1_0_0_R0_MINUS:I I1_1_2_1_0_0_R0_PLUS:I 
*.PININFO I1_1_2_1_1_0_R0_MINUS:I I1_1_2_1_1_0_R0_PLUS:I 
*.PININFO I1_1_2_2_0_0_R0_MINUS:I I1_1_2_2_0_0_R0_PLUS:I 
*.PININFO I1_1_2_2_1_0_R0_MINUS:I I1_1_2_2_1_0_R0_PLUS:I 
*.PININFO I1_2_0_0_0_0_R0_MINUS:I I1_2_0_0_0_0_R0_PLUS:I 
*.PININFO I1_2_0_0_1_0_R0_MINUS:I I1_2_0_0_1_0_R0_PLUS:I 
*.PININFO I1_2_0_1_0_0_R0_MINUS:I I1_2_0_1_0_0_R0_PLUS:I 
*.PININFO I1_2_0_1_1_0_R0_MINUS:I I1_2_0_1_1_0_R0_PLUS:I 
*.PININFO I1_2_0_2_0_0_R0_MINUS:I I1_2_0_2_0_0_R0_PLUS:I 
*.PININFO I1_2_0_2_1_0_R0_MINUS:I I1_2_0_2_1_0_R0_PLUS:I 
*.PININFO I1_2_1_0_0_0_R0_MINUS:I I1_2_1_0_0_0_R0_PLUS:I 
*.PININFO I1_2_1_0_1_0_R0_MINUS:I I1_2_1_0_1_0_R0_PLUS:I 
*.PININFO I1_2_1_1_0_0_R0_MINUS:I I1_2_1_1_0_0_R0_PLUS:I 
*.PININFO I1_2_1_1_1_0_R0_MINUS:I I1_2_1_1_1_0_R0_PLUS:I 
*.PININFO I1_2_1_2_0_0_R0_MINUS:I I1_2_1_2_0_0_R0_PLUS:I 
*.PININFO I1_2_1_2_1_0_R0_MINUS:I I1_2_1_2_1_0_R0_PLUS:I 
*.PININFO I1_2_2_0_0_0_R0_MINUS:I I1_2_2_0_0_0_R0_PLUS:I 
*.PININFO I1_2_2_0_1_0_R0_MINUS:I I1_2_2_0_1_0_R0_PLUS:I 
*.PININFO I1_2_2_1_0_0_R0_MINUS:I I1_2_2_1_0_0_R0_PLUS:I 
*.PININFO I1_2_2_1_1_0_R0_MINUS:I I1_2_2_1_1_0_R0_PLUS:I 
*.PININFO I1_2_2_2_0_0_R0_MINUS:I I1_2_2_2_0_0_R0_PLUS:I 
*.PININFO I1_2_2_2_1_0_R0_MINUS:I I1_2_2_2_1_0_R0_PLUS:I I1_default_MINUS:I 
*.PININFO I1_default_PLUS:I gnd!:I
RI1_2_2_2_1_0_R0 I1_2_2_2_1_0_R0_PLUS I1_2_2_2_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=8.0 l=50u w=50u r=187.206 par=8.0 s=1
RI1_2_2_2_0_0_R0 I1_2_2_2_0_0_R0_PLUS I1_2_2_2_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=50u w=50u r=187.206 par=1.0 s=8
RI1_2_2_1_1_0_R0 I1_2_2_1_1_0_R0_PLUS I1_2_2_1_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=3.0 l=50u w=50u r=187.206 par=3.0 s=1
RI1_2_2_1_0_0_R0 I1_2_2_1_0_0_R0_PLUS I1_2_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=50u w=50u r=187.206 par=1.0 s=3
RI1_2_2_0_1_0_R0 I1_2_2_0_1_0_R0_PLUS I1_2_2_0_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=50u w=50u r=187.206 par=1.0 s=1
RI1_2_2_0_0_0_R0 I1_2_2_0_0_0_R0_PLUS I1_2_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=50u w=50u r=187.206 par=1.0 s=1
RI1_2_1_2_1_0_R0 I1_2_1_2_1_0_R0_PLUS I1_2_1_2_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=8.0 l=7.6u w=50u r=30.1528 par=8.0 s=1
RI1_2_1_2_0_0_R0 I1_2_1_2_0_0_R0_PLUS I1_2_1_2_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=7.6u w=50u r=30.1528 par=1.0 s=8
RI1_2_1_1_1_0_R0 I1_2_1_1_1_0_R0_PLUS I1_2_1_1_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=3.0 l=7.6u w=50u r=30.1528 par=3.0 s=1
RI1_2_1_1_0_0_R0 I1_2_1_1_0_0_R0_PLUS I1_2_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=7.6u w=50u r=30.1528 par=1.0 s=3
RI1_2_1_0_1_0_R0 I1_2_1_0_1_0_R0_PLUS I1_2_1_0_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=7.6u w=50u r=30.1528 par=1.0 s=1
RI1_2_1_0_0_0_R0 I1_2_1_0_0_0_R0_PLUS I1_2_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=7.6u w=50u r=30.1528 par=1.0 s=1
RI1_2_0_2_1_0_R0 I1_2_0_2_1_0_R0_PLUS I1_2_0_2_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=8.0 l=1.6u w=50u r=7.92835 par=8.0 s=1
RI1_2_0_2_0_0_R0 I1_2_0_2_0_0_R0_PLUS I1_2_0_2_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=1.6u w=50u r=7.92835 par=1.0 s=8
RI1_2_0_1_1_0_R0 I1_2_0_1_1_0_R0_PLUS I1_2_0_1_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=3.0 l=1.6u w=50u r=7.92835 par=3.0 s=1
RI1_2_0_1_0_0_R0 I1_2_0_1_0_0_R0_PLUS I1_2_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=1.6u w=50u r=7.92835 par=1.0 s=3
RI1_2_0_0_1_0_R0 I1_2_0_0_1_0_R0_PLUS I1_2_0_0_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=1.6u w=50u r=7.92835 par=1.0 s=1
RI1_2_0_0_0_0_R0 I1_2_0_0_0_0_R0_PLUS I1_2_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=1.6u w=50u r=7.92835 par=1.0 s=1
RI1_1_2_2_1_0_R0 I1_1_2_2_1_0_R0_PLUS I1_1_2_2_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=8.0 l=50u w=3.62u r=2.62272K par=8.0 s=1
RI1_1_2_2_0_0_R0 I1_1_2_2_0_0_R0_PLUS I1_1_2_2_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=50u w=3.62u r=2.62272K par=1.0 s=8
RI1_1_2_1_1_0_R0 I1_1_2_1_1_0_R0_PLUS I1_1_2_1_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=3.0 l=50u w=3.62u r=2.62272K par=3.0 s=1
RI1_1_2_1_0_0_R0 I1_1_2_1_0_0_R0_PLUS I1_1_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=50u w=3.62u r=2.62272K par=1.0 s=3
RI1_1_2_0_1_0_R0 I1_1_2_0_1_0_R0_PLUS I1_1_2_0_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=50u w=3.62u r=2.62272K par=1.0 s=1
RI1_1_2_0_0_0_R0 I1_1_2_0_0_0_R0_PLUS I1_1_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=50u w=3.62u r=2.62272K par=1.0 s=1
RI1_1_1_2_1_0_R0 I1_1_1_2_1_0_R0_PLUS I1_1_1_2_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=8.0 l=7.6u w=3.62u r=422.435 par=8.0 s=1
RI1_1_1_2_0_0_R0 I1_1_1_2_0_0_R0_PLUS I1_1_1_2_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=7.6u w=3.62u r=422.435 par=1.0 s=8
RI1_1_1_1_1_0_R0 I1_1_1_1_1_0_R0_PLUS I1_1_1_1_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=3.0 l=7.6u w=3.62u r=422.435 par=3.0 s=1
RI1_1_1_1_0_0_R0 I1_1_1_1_0_0_R0_PLUS I1_1_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=7.6u w=3.62u r=422.435 par=1.0 s=3
RI1_1_1_0_1_0_R0 I1_1_1_0_1_0_R0_PLUS I1_1_1_0_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=7.6u w=3.62u r=422.435 par=1.0 s=1
RI1_1_1_0_0_0_R0 I1_1_1_0_0_0_R0_PLUS I1_1_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=7.6u w=3.62u r=422.435 par=1.0 s=1
RI1_1_0_2_1_0_R0 I1_1_0_2_1_0_R0_PLUS I1_1_0_2_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=8.0 l=1.6u w=3.62u r=111.075 par=8.0 s=1
RI1_1_0_2_0_0_R0 I1_1_0_2_0_0_R0_PLUS I1_1_0_2_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=1.6u w=3.62u r=111.075 par=1.0 s=8
RI1_1_0_1_1_0_R0 I1_1_0_1_1_0_R0_PLUS I1_1_0_1_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=3.0 l=1.6u w=3.62u r=111.075 par=3.0 s=1
RI1_1_0_1_0_0_R0 I1_1_0_1_0_0_R0_PLUS I1_1_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=1.6u w=3.62u r=111.075 par=1.0 s=3
RI1_1_0_0_1_0_R0 I1_1_0_0_1_0_R0_PLUS I1_1_0_0_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=1.6u w=3.62u r=111.075 par=1.0 s=1
RI1_1_0_0_0_0_R0 I1_1_0_0_0_0_R0_PLUS I1_1_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=1.6u w=3.62u r=111.075 par=1.0 s=1
RI1_0_2_2_1_0_R0 I1_0_2_2_1_0_R0_PLUS I1_0_2_2_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=8.0 l=50u w=800n r=12.5503K par=8.0 s=1
RI1_0_2_2_0_0_R0 I1_0_2_2_0_0_R0_PLUS I1_0_2_2_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=50u w=800n r=12.5503K par=1.0 s=8
RI1_0_2_1_1_0_R0 I1_0_2_1_1_0_R0_PLUS I1_0_2_1_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=3.0 l=50u w=800n r=12.5503K par=3.0 s=1
RI1_0_2_1_0_0_R0 I1_0_2_1_0_0_R0_PLUS I1_0_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=50u w=800n r=12.5503K par=1.0 s=3
RI1_0_2_0_1_0_R0 I1_0_2_0_1_0_R0_PLUS I1_0_2_0_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=50u w=800n r=12.5503K par=1.0 s=1
RI1_0_2_0_0_0_R0 I1_0_2_0_0_0_R0_PLUS I1_0_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=50u w=800n r=12.5503K par=1.0 s=1
RI1_0_1_2_1_0_R0 I1_0_1_2_1_0_R0_PLUS I1_0_1_2_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=8.0 l=7.6u w=800n r=2.02145K par=8.0 s=1
RI1_0_1_2_0_0_R0 I1_0_1_2_0_0_R0_PLUS I1_0_1_2_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=7.6u w=800n r=2.02145K par=1.0 s=8
RI1_0_1_1_1_0_R0 I1_0_1_1_1_0_R0_PLUS I1_0_1_1_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=3.0 l=7.6u w=800n r=2.02145K par=3.0 s=1
RI1_0_1_1_0_0_R0 I1_0_1_1_0_0_R0_PLUS I1_0_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=7.6u w=800n r=2.02145K par=1.0 s=3
RI1_0_1_0_1_0_R0 I1_0_1_0_1_0_R0_PLUS I1_0_1_0_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=7.6u w=800n r=2.02145K par=1.0 s=1
RI1_0_1_0_0_0_R0 I1_0_1_0_0_0_R0_PLUS I1_0_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=7.6u w=800n r=2.02145K par=1.0 s=1
RI1_0_0_2_1_0_R0 I1_0_0_2_1_0_R0_PLUS I1_0_0_2_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=8.0 l=1.6u w=800n r=531.519 par=8.0 s=1
RI1_0_0_2_0_0_R0 I1_0_0_2_0_0_R0_PLUS I1_0_0_2_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=1.6u w=800n r=531.519 par=1.0 s=8
RI1_0_0_1_1_0_R0 I1_0_0_1_1_0_R0_PLUS I1_0_0_1_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=3.0 l=1.6u w=800n r=531.519 par=3.0 s=1
RI1_0_0_1_0_0_R0 I1_0_0_1_0_0_R0_PLUS I1_0_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=1.6u w=800n r=531.519 par=1.0 s=3
RI1_0_0_0_1_0_R0 I1_0_0_0_1_0_R0_PLUS I1_0_0_0_1_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=1.6u w=800n r=531.519 par=1.0 s=1
RI1_0_0_0_0_0_R0 I1_0_0_0_0_0_R0_PLUS I1_0_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[pplus_u] m=1.0 l=1.6u w=800n r=531.519 par=1.0 s=1
RI1_default I1_default_PLUS I1_default_MINUS $SUB=gnd! $[pplus_u] m=1.0 l=2u 
+ w=1u r=497.3349 par=1.0 s=1
.ENDS

