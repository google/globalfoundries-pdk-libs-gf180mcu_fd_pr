* 
* ******************************************************************************
* *                                                                            *
* *                   Copyright 2014, GlobalFoundries                          *
* *                           All rights reserved.                             *
* *                                                                            *
* *                                                                            *
* *                                                                            *
* * This file has been provided pursuant to a License Agreement containing     *
* * restrictions on its use. This file contains valuable trade secrets and     *
* * proprietary information of GlobalFoundries, and is protected by U.S. and   * 
* * international laws and/or treaties.                                        *
* *                                                                            *
* * The copyright notice(s) in this file does not indicate actual or intended  *
* * publication of this file.                                                  *
* *                                                                            *
* * revision: 1.1                                                              *
* ******************************************************************************
* 
* 
* Running on scgtgar01 
* Local time is now Wed, 19 Mar 2014, 11:50:33.
* Main process id is 23919.
*
********************************************************************************
*                                                                              *
* Cellname:   ADDF_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026                                                         *
* at 11:48:26 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************

*.SCALE METER

.SUBCKT ADDF_X1 A B CI CO S VDD VNW VPW VSS 
*.PININFO A:I B:I CI:I CO:O S:O VDD:P VNW:P VPW:P VSS:G 
*.EQN CO=(((B * CI) + (B * A)) + (CI * A));S=!((!((B * CI) + !(B + CI)) * A) + !(!((B * CI) + !(B + CI)) + A))
M_M51 VSS net9 S VPW nmos_5p0 W=1.180000U L=0.600000U
M_M50 net49 A VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_M48 net47 B net49 VPW nmos_5p0 W=0.590000U L=0.600000U
M_M46 net9 CI net47 VPW nmos_5p0 W=0.590000U L=0.600000U
M_M41 net9 net7 net42 VPW nmos_5p0 W=0.590000U L=0.600000U
M_M43 net42 A VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_M44 VSS B net42 VPW nmos_5p0 W=0.590000U L=0.600000U
M_M45 net42 CI VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_M40 VSS B net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_M39 net5 A VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_M38 net7 CI net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_M37 net36 B net7 VPW nmos_5p0 W=0.590000U L=0.600000U
M_M35 VSS A net36 VPW nmos_5p0 W=0.590000U L=0.600000U
M_M34 CO net7 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_M33 VDD net9 S VNW pmos_5p0 W=1.830000U L=0.500000U
M_M32 net31 A VDD VNW pmos_5p0 W=0.990000U L=0.500000U
M_M30 net29 B net31 VNW pmos_5p0 W=0.990000U L=0.500000U
M_M28 net9 CI net29 VNW pmos_5p0 W=0.990000U L=0.500000U
M_M24 net9 net7 net3 VNW pmos_5p0 W=0.990000U L=0.500000U
M_M25 net3 A VDD VNW pmos_5p0 W=0.990000U L=0.500000U
M_M26 VDD B net3 VNW pmos_5p0 W=0.990000U L=0.500000U
M_M27 net3 CI VDD VNW pmos_5p0 W=0.990000U L=0.500000U
M_M23 VDD B net1 VNW pmos_5p0 W=0.990000U L=0.500000U
M_M22 net1 A VDD VNW pmos_5p0 W=0.990000U L=0.500000U
M_M21 net7 CI net1 VNW pmos_5p0 W=0.990000U L=0.500000U
M_M20 net19 B net7 VNW pmos_5p0 W=0.990000U L=0.500000U
M_M18 VDD A net19 VNW pmos_5p0 W=0.990000U L=0.500000U
M_M17 CO net7 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   ADDF_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:48:24 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT ADDF_X2 A B CI CO S VDD VNW VPW VSS 
*.PININFO A:I B:I CI:I CO:O S:O VDD:P VNW:P VPW:P VSS:G 
*.EQN CO=(((B * CI) + (B * A)) + (CI * A));S=!((!((B * CI) + !(B + CI)) * A) + !(!((B * CI) + !(B + CI)) + A))
M_M51_17 VSS net9 S VPW nmos_5p0 W=1.320000U L=0.600000U
M_M51 VSS net9 S VPW nmos_5p0 W=1.320000U L=0.600000U
M_M50 net49 A VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_M48 net47 B net49 VPW nmos_5p0 W=0.800000U L=0.600000U
M_M46 net9 CI net47 VPW nmos_5p0 W=0.800000U L=0.600000U
M_M41 net9 net7 net42 VPW nmos_5p0 W=0.800000U L=0.600000U
M_M43 net42 A VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_M44 VSS B net42 VPW nmos_5p0 W=0.800000U L=0.600000U
M_M45 net42 CI VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_M40 VSS B net5 VPW nmos_5p0 W=0.800000U L=0.600000U
M_M39 net5 A VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_M38 net7 CI net5 VPW nmos_5p0 W=0.800000U L=0.600000U
M_M37 net36 B net7 VPW nmos_5p0 W=0.800000U L=0.600000U
M_M35 VSS A net36 VPW nmos_5p0 W=0.800000U L=0.600000U
M_M34 CO net7 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_M34_25 CO net7 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_M33_12 VDD net9 S VNW pmos_5p0 W=1.800000U L=0.500000U
M_M33 VDD net9 S VNW pmos_5p0 W=1.800000U L=0.500000U
M_M32 net31 A VDD VNW pmos_5p0 W=1.390000U L=0.500000U
M_M30 net29 B net31 VNW pmos_5p0 W=1.390000U L=0.500000U
M_M28 net9 CI net29 VNW pmos_5p0 W=1.390000U L=0.500000U
M_M24 net9 net7 net3 VNW pmos_5p0 W=1.390000U L=0.500000U
M_M25 net3 A VDD VNW pmos_5p0 W=1.390000U L=0.500000U
M_M26 VDD B net3 VNW pmos_5p0 W=1.390000U L=0.500000U
M_M27 net3 CI VDD VNW pmos_5p0 W=1.390000U L=0.500000U
M_M23 VDD B net1 VNW pmos_5p0 W=1.390000U L=0.500000U
M_M22 net1 A VDD VNW pmos_5p0 W=1.390000U L=0.500000U
M_M21 net7 CI net1 VNW pmos_5p0 W=1.390000U L=0.500000U
M_M20 net19 B net7 VNW pmos_5p0 W=1.390000U L=0.500000U
M_M18 VDD A net19 VNW pmos_5p0 W=1.390000U L=0.500000U
M_M17 CO net7 VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_M17_23 CO net7 VDD VNW pmos_5p0 W=1.800000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   ADDF_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs008             *
* at 11:48:24 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT ADDF_X4 A B CI CO S VDD VNW VPW VSS 
*.PININFO A:I B:I CI:I CO:O S:O VDD:P VNW:P VPW:P VSS:G 
*.EQN CO=(((B * CI) + (B * A)) + (CI * A));S=!((!((B * CI) + !(B + CI)) * A) + !(!((B * CI) + !(B + CI)) + A))
M_M51_17_0 VSS net9 S VPW nmos_5p0 W=1.320000U L=0.600000U
M_M51_18 VSS net9 S VPW nmos_5p0 W=1.320000U L=0.600000U
M_M51_17 VSS net9 S VPW nmos_5p0 W=1.320000U L=0.600000U
M_M51 VSS net9 S VPW nmos_5p0 W=1.320000U L=0.600000U
M_M50 net49 A VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_M48 net47 B net49 VPW nmos_5p0 W=0.800000U L=0.600000U
M_M46 net9 CI net47 VPW nmos_5p0 W=0.800000U L=0.600000U
M_M41 net9 net7 net42 VPW nmos_5p0 W=0.800000U L=0.600000U
M_M43 net42 A VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_M44 VSS B net42 VPW nmos_5p0 W=0.800000U L=0.600000U
M_M45 net42 CI VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_M40 VSS B net5 VPW nmos_5p0 W=0.800000U L=0.600000U
M_M39 net5 A VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_M38 net7 CI net5 VPW nmos_5p0 W=0.800000U L=0.600000U
M_M37 net36 B net7 VPW nmos_5p0 W=0.800000U L=0.600000U
M_M35 VSS A net36 VPW nmos_5p0 W=0.800000U L=0.600000U
M_M34 CO net7 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_M34_25 CO net7 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_M34_53 CO net7 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_M34_25_56 CO net7 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_M33_12_23 VDD net9 S VNW pmos_5p0 W=1.830000U L=0.500000U
M_M33_34 VDD net9 S VNW pmos_5p0 W=1.830000U L=0.500000U
M_M33_12 VDD net9 S VNW pmos_5p0 W=1.830000U L=0.500000U
M_M33 VDD net9 S VNW pmos_5p0 W=1.830000U L=0.500000U
M_M32 net31 A VDD VNW pmos_5p0 W=1.390000U L=0.500000U
M_M30 net29 B net31 VNW pmos_5p0 W=1.390000U L=0.500000U
M_M28 net9 CI net29 VNW pmos_5p0 W=1.390000U L=0.500000U
M_M24 net9 net7 net3 VNW pmos_5p0 W=1.390000U L=0.500000U
M_M25 net3 A VDD VNW pmos_5p0 W=1.390000U L=0.500000U
M_M26 VDD B net3 VNW pmos_5p0 W=1.390000U L=0.500000U
M_M27 net3 CI VDD VNW pmos_5p0 W=1.390000U L=0.500000U
M_M23 VDD B net1 VNW pmos_5p0 W=1.390000U L=0.500000U
M_M22 net1 A VDD VNW pmos_5p0 W=1.390000U L=0.500000U
M_M21 net7 CI net1 VNW pmos_5p0 W=1.390000U L=0.500000U
M_M20 net19 B net7 VNW pmos_5p0 W=1.390000U L=0.500000U
M_M18 VDD A net19 VNW pmos_5p0 W=1.390000U L=0.500000U
M_M17 CO net7 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_M17_23 CO net7 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_M17_66 CO net7 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_M17_23_46 CO net7 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   ADDH_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:42 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT ADDH_X1 A B CO S VDD VNW VPW VSS 
*.PININFO A:I B:I CO:O S:O VDD:P VNW:P VPW:P VSS:G 
*.EQN CO=(A * B);S=!((A * B) + !(A + B))
M_i_2 VSS NCO CO VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5 net_0 A VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_4 NCO B net_0 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_9 NS B net_1 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_8 net_1 A NS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_10 VSS NCO net_1 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_0 S NS VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 VDD NCO CO VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7 NCO A VDD VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_6 VDD B NCO VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_12 net_2 B VDD VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_11 NS A net_2 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_13 VDD NCO NS VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_1 S NS VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   ADDH_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:48:37 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT ADDH_X2 A B CO S VDD VNW VPW VSS 
*.PININFO A:I B:I CO:O S:O VDD:P VNW:P VPW:P VSS:G 
*.EQN CO=(A * B);S=!((A * B) + !(A + B))
M_i_2_1 CO NCO VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 VSS NCO CO VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5 net_0 A VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4 NCO B net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_9 NS B net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_8 net_1 A NS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_10 VSS NCO net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 S NS VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 VSS NS S VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 CO NCO VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0 VDD NCO CO VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7 NCO A VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 VDD B NCO VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_12 net_2 B VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11 NS A net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_13 VDD NCO NS VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 S NS VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 VDD NS S VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   ADDH_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:44 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT ADDH_X4 A B CO S VDD VNW VPW VSS 
*.PININFO A:I B:I CO:O S:O VDD:P VNW:P VPW:P VSS:G 
*.EQN CO=(A * B);S=!((A * B) + !(A + B))
M_i_5_1 net_0_0 A VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_1 NCO B net_0_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_0 net_0_1 B NCO VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_0 VSS A net_0_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_10_0 net_1 NCO VSS VPW nmos_5p0 W=0.880000U L=0.600000U
M_i_8_0 NS A net_1 VPW nmos_5p0 W=0.880000U L=0.600000U
M_i_9_0 net_1 B NS VPW nmos_5p0 W=0.880000U L=0.600000U
M_i_9_1 NS B net_1 VPW nmos_5p0 W=0.880000U L=0.600000U
M_i_8_1 net_1 A NS VPW nmos_5p0 W=0.880000U L=0.600000U
M_i_10_1 VSS NCO net_1 VPW nmos_5p0 W=0.880000U L=0.600000U
M_i_2_3 CO NCO VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_2 VSS NCO CO VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 CO NCO VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 VSS NCO CO VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 S NS VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 VSS NS S VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 S NS VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 VSS NS S VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_7_1 NCO A VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 VDD B NCO VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 NCO B VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 VDD A NCO VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_13_0 NS NCO VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_0 net_2_0 A NS VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_12_0 VDD B net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_12_1 net_2_1 B VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_1 NS A net_2_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_13_1 VDD NCO NS VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_3 CO NCO VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_2 VDD NCO CO VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 CO NCO VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0 VDD NCO CO VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 S NS VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 VDD NS S VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 S NS VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 VDD NS S VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AND2_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:36 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AND2_X1 A1 A2 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=(A1 * A2)
M_i_2 net_0 A1 Z_neg VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_3 VSS A2 net_0 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4 Z_neg A1 VDD VNW pmos_5p0 W=0.820000U L=0.500000U
M_i_5 VDD A2 Z_neg VNW pmos_5p0 W=0.820000U L=0.500000U
M_i_1 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AND2_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:48:35 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AND2_X2 A1 A2 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=(A1 * A2)
M_i_2 net_0 A1 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 VSS A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4 Z_neg A1 VDD VNW pmos_5p0 W=1.640000U L=0.500000U
M_i_5 VDD A2 Z_neg VNW pmos_5p0 W=1.640000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AND2_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:48:35 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AND2_X4 A1 A2 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=(A1 * A2)
M_i_3_1 net_0_1 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 Z_neg A1 net_0_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_0_0 A1 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 VSS A2 net_0_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_1 Z_neg A2 VDD VNW pmos_5p0 W=1.640000U L=0.500000U
M_i_4_1 VDD A1 Z_neg VNW pmos_5p0 W=1.640000U L=0.500000U
M_i_4_0 Z_neg A1 VDD VNW pmos_5p0 W=1.640000U L=0.500000U
M_i_5_0 VDD A2 Z_neg VNW pmos_5p0 W=1.640000U L=0.500000U
M_i_1_3 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AND3_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs024             *
* at 11:48:19 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AND3_X1 A1 A2 A3 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=((A1 * A2) * A3)
M_i_2 net_0 A1 Z_neg VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_3 net_1 A2 net_0 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_4 VSS A3 net_1 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5 VDD A1 Z_neg VNW pmos_5p0 W=0.730000U L=0.500000U
M_i_6 Z_neg A2 VDD VNW pmos_5p0 W=0.730000U L=0.500000U
M_i_7 VDD A3 Z_neg VNW pmos_5p0 W=0.730000U L=0.500000U
M_i_1 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AND3_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs008             *
* at 11:48:15 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AND3_X2 A1 A2 A3 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=((A1 * A2) * A3)
M_i_2 net_0 A1 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 net_1 A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4 VSS A3 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5 VDD A1 Z_neg VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_6 Z_neg A2 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_7 VDD A3 Z_neg VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AND3_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs027             *
* at 11:48:16 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AND3_X4 A1 A2 A3 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=((A1 * A2) * A3)
M_i_4_0 net_1_1 A3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 net_0_1 A2 net_1_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 Z_neg A1 net_0_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_0_0 A1 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 net_1_0 A2 net_0_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_1 VSS A3 net_1_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_7_0 Z_neg A3 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_6_1 VDD A2 Z_neg VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_5_1 Z_neg A1 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_5_0 VDD A1 Z_neg VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_6_0 Z_neg A2 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_7_1 VDD A3 Z_neg VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_1_3 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AND4_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:02 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AND4_X1 A1 A2 A3 A4 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I A4:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=(((A1 * A2) * A3) * A4)
M_i_2 net_0 A1 Z_neg VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_3 net_1 A2 net_0 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_4 net_2 A3 net_1 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_5 VSS A4 net_2 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6 Z_neg A1 VDD VNW pmos_5p0 W=0.640000U L=0.500000U
M_i_7 VDD A2 Z_neg VNW pmos_5p0 W=0.640000U L=0.500000U
M_i_8 Z_neg A3 VDD VNW pmos_5p0 W=0.640000U L=0.500000U
M_i_9 VDD A4 Z_neg VNW pmos_5p0 W=0.640000U L=0.500000U
M_i_1 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AND4_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:04 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AND4_X2 A1 A2 A3 A4 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I A4:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=(((A1 * A2) * A3) * A4)
M_i_2 net_0 A1 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 net_1 A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4 net_2 A3 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5 VSS A4 net_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6 Z_neg A1 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_7 VDD A2 Z_neg VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_8 Z_neg A3 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_9 VDD A4 Z_neg VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AND4_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:04 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AND4_X4 A1 A2 A3 A4 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I A4:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=(((A1 * A2) * A3) * A4)
M_i_5_1 net_2_1 A4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_1 net_1_1 A3 net_2_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 net_0_1 A2 net_1_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 Z_neg A1 net_0_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_0_0 A1 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 net_1_0 A2 net_0_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_0 net_2_0 A3 net_1_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_0 VSS A4 net_2_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_9_1 Z_neg A4 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_8_1 VDD A3 Z_neg VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_7_1 Z_neg A2 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_6_1 VDD A1 Z_neg VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_6_0 Z_neg A1 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_7_0 VDD A2 Z_neg VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_8_0 Z_neg A3 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_9_0 VDD A4 Z_neg VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_1_3 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI211_X1.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:01 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AOI211_X1 A1 A2 B C ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B:I C:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 * A2) + B) + C)
M_i_1 net_0 A2 VSS VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_0 ZN A1 net_0 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_2 VSS B ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_3 ZN C VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_5 ZN A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4 net_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 net_2 B net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7 VDD C net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI211_X2.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:02 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AOI211_X2 A1 A2 B C ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B:I C:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 * A2) + B) + C)
M_i_1_1 net_0_0 A2 VSS VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_0_1 ZN A1 net_0_0 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_0_0 net_0_1 A1 ZN VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_1_0 VSS A2 net_0_1 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_2_0 ZN B VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_3_0 VSS C ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_3_1 ZN C VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_2_1 VSS B ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_5_1 ZN A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 net_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 ZN A1 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 net_1 A2 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 net_2_0 B net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 VDD C net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 net_2_1 C VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 net_1 B net_2_1 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI211_X4.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:06 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AOI211_X4 A1 A2 B C ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B:I C:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 * A2) + B) + C)
M_i_1_3 net_0_0 A2 VSS VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_0_3 ZN A1 net_0_0 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_0_2 net_0_1 A1 ZN VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_1_2 VSS A2 net_0_1 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_1_1 net_0_2 A2 VSS VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_0_1 ZN A1 net_0_2 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_0_0 net_0_3 A1 ZN VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_1_0 VSS A2 net_0_3 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_2_0 ZN B VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_3_0 VSS C ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_3_1 ZN C VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_2_1 VSS B ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_2_2 ZN B VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_3_2 VSS C ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_3_3 ZN C VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_2_3 VSS B ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_5_3 ZN A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_3 net_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_2 ZN A1 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_2 net_1 A2 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 ZN A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 net_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 ZN A1 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 net_1 A2 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 net_2_0 B net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 VDD C net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 net_2_1 C VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 net_1 B net_2_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_2 net_2_2 B net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_2 VDD C net_2_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_3 net_2_3 C VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_3 net_1 B net_2_3 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI21_X1.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:48:13 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AOI21_X1 A1 A2 B ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!((A1 * A2) + B)
M_i_1 net_0 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2 VSS B ZN VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_4 ZN A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3 net_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5 VDD B net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI21_X2.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs007             *
* at 11:48:13 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AOI21_X2 A1 A2 B ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!((A1 * A2) + B)
M_i_2_0 ZN B VSS VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_2_1 VSS B ZN VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_1_0 net_0_0 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 ZN A1 net_0_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 net_0_1 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 VSS A2 net_0_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_0 VDD B net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 net_1 B VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 ZN A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 net_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0 ZN A1 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 net_1 A2 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI21_X4.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs007             *
* at 11:48:12 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AOI21_X4 A1 A2 B ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!((A1 * A2) + B)
M_i_1_3 net_0_0 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 ZN A1 net_0_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 net_0_1 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_2 VSS A2 net_0_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 net_0_2 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 ZN A1 net_0_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 net_0_3 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 VSS A2 net_0_3 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_3 ZN B VSS VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_2_2 VSS B ZN VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_2_1 ZN B VSS VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_2_0 VSS B ZN VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_4_3 ZN A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_3 net_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_2 ZN A1 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_2 net_1 A2 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 ZN A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 net_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0 ZN A1 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 net_1 A2 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_3 VDD B net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_2 net_1 B VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 VDD B net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 net_1 B VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI221_X1.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:47:43 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AOI221_X1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B1:I B2:I C:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 * A2) + (B1 * B2)) + C)
M_i_4 net_1 B2 VSS VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_3 ZN B1 net_1 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_2 VSS C ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_1 net_0 A2 VSS VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_0 ZN A1 net_0 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_9 VDD B2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8 net_3 B1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7 net_2 C net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 ZN A2 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5 net_2 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI221_X2.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs010             *
* at 11:47:44 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AOI221_X2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B1:I B2:I C:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 * A2) + (B1 * B2)) + C)
M_i_2_1 VSS C ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_4_1 net_1_0 B2 VSS VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_3_1 ZN B1 net_1_0 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_3_0 net_1_1 B1 ZN VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_4_0 VSS B2 net_1_1 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_2_0 ZN C VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_0_1 net_0_0 A1 ZN VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_1_1 VSS A2 net_0_0 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_1_0 net_0_1 A2 VSS VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_0_0 ZN A1 net_0_1 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_7_1 net_3 C net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_1 VDD B2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_1 net_3 B1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_0 VDD B1 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_0 net_3 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 net_2 C net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 ZN A1 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 net_2 A2 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 ZN A2 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 net_2 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI221_X4.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:47:50 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AOI221_X4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B1:I B2:I C:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 * A2) + (B1 * B2)) + C)
M_i_3_3 net_1_0 B1 ZN VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_4_3 VSS B2 net_1_0 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_4_2 net_1_1 B2 VSS VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_3_2 ZN B1 net_1_1 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_3_1 net_1_2 B1 ZN VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_4_1 VSS B2 net_1_2 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_4_0 net_1_3 B2 VSS VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_3_0 ZN B1 net_1_3 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_2_3 VSS C ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_2_2 ZN C VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_2_1 VSS C ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_2_0 ZN C VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_0_3 net_0_0 A1 ZN VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_1_3 VSS A2 net_0_0 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_1_2 net_0_1 A2 VSS VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_0_2 ZN A1 net_0_1 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_0_1 net_0_2 A1 ZN VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_1_1 VSS A2 net_0_2 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_1_0 net_0_3 A2 VSS VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_0_0 ZN A1 net_0_3 VPW nmos_5p0 W=1.185000U L=0.600000U
M_i_8_3 net_3 B1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_3 VDD B2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_2 net_3 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_2 VDD B1 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_1 net_3 B1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_1 VDD B2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_0 net_3 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_0 VDD B1 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_3 net_3 C net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_2 net_2 C net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 net_3 C net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 net_2 C net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_3 ZN A1 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_3 net_2 A2 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_2 ZN A2 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_2 net_2 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 ZN A1 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 net_2 A2 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 ZN A2 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 net_2 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI222_X1.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:47:39 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AOI222_X1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 * A2) + (B1 * B2)) + (C1 * C2))
M_i_5 net_2 C2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4 ZN C1 net_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2 net_1 B1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 VSS B2 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1 net_0 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_11 net_4 C2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10 VDD C1 net_4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8 net_4 B1 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9 net_3 B2 net_4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7 ZN A2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 net_3 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI222_X2.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:47:41 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AOI222_X2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 * A2) + (B1 * B2)) + (C1 * C2))
M_i_4_1 net_2_1 C1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_1 VSS C2 net_2_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_0 net_2_0 C2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_0 ZN C1 net_2_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_1_1 B1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 VSS B2 net_1_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 net_1_0 B2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 ZN B1 net_1_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 net_0_1 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 VSS A2 net_0_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 net_0_0 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 ZN A1 net_0_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_10_1 net_4 C1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_1 VDD C2 net_4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_0 net_4 C2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10_0 VDD C1 net_4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_0 net_4 B1 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_0 net_3 B2 net_4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_1 net_4 B2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_1 net_3 B1 net_4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 ZN A1 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 net_3 A2 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 ZN A2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 net_3 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI222_X4.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:47:44 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AOI222_X4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 * A2) + (B1 * B2)) + (C1 * C2))
M_i_4_3 net_2_3 C1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_3 VSS C2 net_2_3 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_2 net_2_2 C2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_2 ZN C1 net_2_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_1 net_2_1 C1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_1 VSS C2 net_2_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_0 net_2_0 C2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_0 ZN C1 net_2_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_1_3 B1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 VSS B2 net_1_3 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 net_1_2 B2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 ZN B1 net_1_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_2 net_1_1 B1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_2 VSS B2 net_1_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_3 net_1_0 B2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_3 ZN B1 net_1_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 net_0_3 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 VSS A2 net_0_3 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 net_0_2 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 ZN A1 net_0_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 net_0_1 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_2 VSS A2 net_0_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_3 net_0_0 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 ZN A1 net_0_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_10_3 net_4 C1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_3 VDD C2 net_4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_2 net_4 C2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10_2 VDD C1 net_4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10_1 net_4 C1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_1 VDD C2 net_4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_0 net_4 C2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10_0 VDD C1 net_4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_0 net_4 B1 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_0 net_3 B2 net_4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_1 net_4 B2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_1 net_3 B1 net_4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_2 net_4 B1 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_2 net_3 B2 net_4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_3 net_4 B2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_3 net_3 B1 net_4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 ZN A1 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 net_3 A2 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 ZN A2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 net_3 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_2 ZN A1 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_2 net_3 A2 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_3 ZN A2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_3 net_3 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI22_X1.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:02 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AOI22_X1 A1 A2 B1 B2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B1:I B2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!((A1 * A2) + (B1 * B2))
M_i_3 net_1 B2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2 ZN B1 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1 VSS A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_7 VDD B2 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 net_2 B1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4 ZN A1 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5 net_2 A2 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI22_X2.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:48:03 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AOI22_X2 A1 A2 B1 B2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B1:I B2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!((A1 * A2) + (B1 * B2))
M_i_3_1 net_1_0 B2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 ZN B1 net_1_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_1_1 B1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 VSS B2 net_1_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 net_0_0 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 ZN A1 net_0_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 net_0_1 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 VSS A2 net_0_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_7_1 VDD B2 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 net_2 B1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 VDD B1 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 net_2 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 ZN A2 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 net_2 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 ZN A1 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 net_2 A2 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   AOI22_X4.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:07 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT AOI22_X4 A1 A2 B1 B2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B1:I B2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!((A1 * A2) + (B1 * B2))
M_i_3_3 net_1_0 B2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_3 ZN B1 net_1_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_2 net_1_1 B1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_2 VSS B2 net_1_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 net_1_2 B2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 ZN B1 net_1_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_1_3 B1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 VSS B2 net_1_3 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 net_0_0 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 ZN A1 net_0_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 net_0_1 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 VSS A2 net_0_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_2 net_0_2 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 ZN A1 net_0_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 net_0_3 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_3 VSS A2 net_0_3 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_7_3 VDD B2 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_3 net_2 B1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_2 VDD B1 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_2 net_2 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 VDD B2 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 net_2 B1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 VDD B1 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 net_2 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 ZN A2 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 net_2 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 ZN A1 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 net_2 A2 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_2 ZN A2 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_2 net_2 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_3 ZN A1 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_3 net_2 A2 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUFZ_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:34 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT BUFZ_X1 EN I Z VDD VNW VPW VSS 
*.PININFO EN:I I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_XX27 VSS EN NEN VPW nmos_5p0 W=0.590000U L=0.600000U
M_XX44 VSS NEN NI_N VPW nmos_5p0 W=0.590000U L=0.600000U
M_XX36 NI_N EN NI_P VPW nmos_5p0 W=0.590000U L=0.600000U
M_XX43 NI_N I VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_XX22 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX28 VDD EN NEN VNW pmos_5p0 W=0.990000U L=0.500000U
M_XX45 NI_P EN VDD VNW pmos_5p0 W=0.990000U L=0.500000U
M_XX39 NI_N NEN NI_P VNW pmos_5p0 W=0.990000U L=0.500000U
M_XX46 NI_P I VDD VNW pmos_5p0 W=0.990000U L=0.500000U
M_XX21 VDD NI_P Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUFZ_X12.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:48:43 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT BUFZ_X12 EN I Z VDD VNW VPW VSS 
*.PININFO EN:I I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_mn VSS EN NEN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn8 NI_N NEN VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn21 NI_P EN NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17 NI_N I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9 VSS I NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_10 NI_N I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9_17 VSS I NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_10_0 NI_N I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9_17_30 VSS I NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25_34 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49_88 VSS NI_N Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_33 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_99 VSS NI_N Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49 VSS NI_N Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3 VSS NI_N Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25_35 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49_80 VSS NI_N Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_34 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_89 VSS NI_N Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_mp VDD EN NEN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp7 NI_P EN VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp22 NI_N NEN NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14 NI_P I VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10 VDD I NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_11 NI_P I VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10_8 VDD I NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_11_21 NI_P I VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10_8_17 VDD I NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57_75 Z NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56_111 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_106 Z NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_58 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57 Z NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12 Z NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57_69 Z NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56_105 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_96 Z NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_57 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUFZ_X16.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:48:47 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT BUFZ_X16 EN I Z VDD VNW VPW VSS 
*.PININFO EN:I I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_mn VSS EN NEN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn8 NI_N NEN VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn21 NI_P EN NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17 NI_N I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9 VSS I NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_10 NI_N I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9_17 VSS I NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_34 NI_N I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9_41 VSS I NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_10_30 NI_N I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9_17_61 VSS I NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25_34 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49_88 VSS NI_N Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_33 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_99 VSS NI_N Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49 VSS NI_N Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3 VSS NI_N Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25_34_75 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49_88_82 VSS NI_N Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_33_198 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_99_125 VSS NI_N Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25_137 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49_181 VSS NI_N Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_65 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_118 VSS NI_N Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_mp VDD EN NEN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp7 NI_P EN VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp22 NI_N NEN NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14 NI_P I VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10 VDD I NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_11 NI_P I VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10_8 VDD I NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_7 NI_P I VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10_32 VDD I NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_11_55 NI_P I VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10_8_20 VDD I NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57_75 Z NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56_111 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_106 Z NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_58 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57 Z NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12 Z NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57_75_85 Z NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56_111_134 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_106_111 Z NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_58_95 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57_97 Z NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56_133 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_126 Z NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_153 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUFZ_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs008             *
* at 11:48:33 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT BUFZ_X2 EN I Z VDD VNW VPW VSS 
*.PININFO EN:I I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_XX27 VSS EN NEN VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX44 VSS NEN NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX36 NI_N EN NI_P VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX43 NI_N I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX22 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX22_4 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX28 VDD EN NEN VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX45 NI_P EN VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX39 NI_N NEN NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX46 NI_P I VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX21 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX21_5 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUFZ_X3.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs010             *
* at 11:48:34 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT BUFZ_X3 EN I Z VDD VNW VPW VSS 
*.PININFO EN:I I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_XX27 VSS EN NEN VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX44 VSS NEN NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX36 NI_N EN NI_P VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX43 NI_N I VSS VPW nmos_5p0 W=0.885000U L=0.600000U
M_XX43_17 NI_N I VSS VPW nmos_5p0 W=0.885000U L=0.600000U
M_XX22 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX22_4 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX22_4_97 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX28 VDD EN NEN VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX45 NI_P EN VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX39 NI_N NEN NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX46 NI_P I VDD VNW pmos_5p0 W=1.485000U L=0.500000U
M_XX46_9 NI_P I VDD VNW pmos_5p0 W=1.485000U L=0.500000U
M_XX21 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX21_5 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX21_5_72 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUFZ_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:48:34 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT BUFZ_X4 EN I Z VDD VNW VPW VSS 
*.PININFO EN:I I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_XX27 VSS EN NEN VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX44 VSS NEN NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX36 NI_N EN NI_P VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX43 NI_N I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX43_17 NI_N I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX22 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX22_4 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX22_4_97 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX22_4_97_16 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX28 VDD EN NEN VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX45 NI_P EN VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX39 NI_N NEN NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX46 NI_P I VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX46_9 NI_P I VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX21 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX21_5 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX21_5_72 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX21_5_72_5 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUFZ_X8.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:48:38 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT BUFZ_X8 EN I Z VDD VNW VPW VSS 
*.PININFO EN:I I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_mn VSS EN NEN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn8 NI_N NEN VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn21 NI_P EN NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17 NI_N I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9 VSS I NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_10 NI_N I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9_17 VSS I NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25_34 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49_88 VSS NI_N Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_33 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_99 VSS NI_N Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49 VSS NI_N Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3 VSS NI_N Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_mp VDD EN NEN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp7 NI_P EN VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp22 NI_N NEN NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14 NI_P I VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10 VDD I NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_11 NI_P I VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10_8 VDD I NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57_75 Z NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56_111 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_106 Z NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_58 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57 Z NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12 Z NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4 VDD NI_P Z VNW pmos_5p0 W=1.800000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUF_X1.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs008             *
* at 11:48:56 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT BUF_X1 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2 VSS I Z_neg VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 VDD I Z_neg VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_1 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUF_X12.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:49:03 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT BUF_X12 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 VSS I Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_2 Z_neg I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_3 VSS I Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_4 Z_neg I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_5 VSS I Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_4 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_5 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_6 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_7 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_8 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_9 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_10 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_11 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_2 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_3 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_4 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_5 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_4 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_5 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_6 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_7 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_8 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_9 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_10 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_11 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUF_X16.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:49:03 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT BUF_X16 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 VSS I Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_2 Z_neg I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_3 VSS I Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_4 Z_neg I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_5 VSS I Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_6 Z_neg I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_7 VSS I Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_4 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_5 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_6 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_7 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_8 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_9 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_10 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_11 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_12 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_13 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_14 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_15 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_2 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_3 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_4 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_5 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_6 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_7 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_4 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_5 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_6 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_7 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_8 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_9 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_10 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_11 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_12 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_13 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_14 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_15 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUF_X2.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs007             *
* at 11:48:56 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT BUF_X2 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2 VSS I Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUF_X20.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:49:10 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT BUF_X20 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 VSS I Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_2 Z_neg I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_3 VSS I Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_4 Z_neg I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_5 VSS I Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_6 Z_neg I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_7 VSS I Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_8 Z_neg I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_9 VSS I Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_4 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_5 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_6 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_7 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_8 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_9 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_10 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_11 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_12 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_13 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_14 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_15 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_16 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_17 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_18 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_19 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_2 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_3 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_4 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_5 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_6 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_7 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_8 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_9 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_4 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_5 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_6 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_7 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_8 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_9 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_10 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_11 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_12 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_13 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_14 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_15 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_16 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_17 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_18 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_19 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUF_X3.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:48:57 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT BUF_X3 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2 VSS I Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUF_X4.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:48:53 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT BUF_X4 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 VSS I Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   BUF_X8.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs010             *
* at 11:48:54 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT BUF_X8 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 VSS I Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_2 Z_neg I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_3 VSS I Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_4 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_5 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_6 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_7 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_2 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_3 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_4 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_5 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_6 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_7 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKBUF_X1.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:48:51 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT CLKBUF_X1 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2 VSS I Z_neg VPW nmos_5p0 W=0.365000U L=0.600000U
M_i_0 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_3 VDD I Z_neg VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_1 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKBUF_X12.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs024             *
* at 11:48:58 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT CLKBUF_X12 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_1 VSS I Z_neg VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_2 Z_neg I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_3 VSS I Z_neg VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_4 Z_neg I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_5 VSS I Z_neg VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_2 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_3 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_4 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_5 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_6 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_7 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_8 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_9 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_10 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_11 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_2 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_3 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_4 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_5 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_4 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_5 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_6 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_7 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_8 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_9 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_10 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_11 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKBUF_X16.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs008             *
* at 11:48:56 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT CLKBUF_X16 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_1 VSS I Z_neg VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_2 Z_neg I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_3 VSS I Z_neg VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_4 Z_neg I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_5 VSS I Z_neg VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_6 Z_neg I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_7 VSS I Z_neg VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_2 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_3 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_4 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_5 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_6 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_7 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_8 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_9 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_10 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_11 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_12 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_13 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_14 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_15 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_2 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_3 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_4 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_5 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_6 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_7 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_4 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_5 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_6 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_7 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_8 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_9 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_10 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_11 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_12 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_13 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_14 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_15 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKBUF_X2.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:48:50 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT CLKBUF_X2 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2 VSS I Z_neg VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_3 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKBUF_X20.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:49:08 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT CLKBUF_X20 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_1 VSS I Z_neg VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_2 Z_neg I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_3 VSS I Z_neg VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_4 Z_neg I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_5 VSS I Z_neg VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_6 Z_neg I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_7 VSS I Z_neg VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_8 Z_neg I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_9 VSS I Z_neg VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_2 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_3 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_4 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_5 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_6 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_7 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_8 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_9 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_10 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_11 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_12 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_13 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_14 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_15 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_16 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_17 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_18 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_19 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_2 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_3 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_4 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_5 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_6 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_7 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_8 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_9 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_4 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_5 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_6 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_7 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_8 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_9 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_10 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_11 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_12 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_13 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_14 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_15 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_16 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_17 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_18 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_19 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKBUF_X3.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs021             *
* at 11:48:53 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT CLKBUF_X3 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.550000U L=0.600000U
M_i_2_1 VSS I Z_neg VPW nmos_5p0 W=0.550000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=0.600000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=0.600000U L=0.600000U
M_i_0_2 Z Z_neg VSS VPW nmos_5p0 W=0.600000U L=0.600000U
M_i_0_3 VSS Z_neg Z VPW nmos_5p0 W=0.600000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=1.375000U L=0.500000U
M_i_3_1 VDD I Z_neg VNW pmos_5p0 W=1.375000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.375000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.375000U L=0.500000U
M_i_1_2 Z Z_neg VDD VNW pmos_5p0 W=1.375000U L=0.500000U
M_i_1_3 VDD Z_neg Z VNW pmos_5p0 W=1.375000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKBUF_X4.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:48:53 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT CLKBUF_X4 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_1 VSS I Z_neg VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_2 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_3 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKBUF_X8.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:56 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT CLKBUF_X8 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_1 VSS I Z_neg VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_2 Z_neg I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_2_3 VSS I Z_neg VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_2 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_3 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_4 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_5 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_6 Z Z_neg VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_0_7 VSS Z_neg Z VPW nmos_5p0 W=0.800000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_2 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_3 VDD I Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_4 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_5 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_6 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_7 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKINV_X1.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs007             *
* at 11:48:46 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT CLKINV_X1 I ZN VDD VNW VPW VSS 
*.PININFO I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_i_0 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_1 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKINV_X12.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:48 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT CLKINV_X12 I ZN VDD VNW VPW VSS 
*.PININFO I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_i_0_0 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_1 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_2 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_3 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_4 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_5 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_6 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_7 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_8 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_9 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_10 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_11 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_1_0 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_4 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_5 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_6 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_7 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_8 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_9 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_10 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_11 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKINV_X16.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:48:50 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT CLKINV_X16 I ZN VDD VNW VPW VSS 
*.PININFO I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_i_0_0 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_1 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_2 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_3 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_4 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_5 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_6 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_7 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_8 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_9 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_10 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_11 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_12 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_13 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_14 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_15 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_1_0 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_4 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_5 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_6 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_7 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_8 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_9 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_10 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_11 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_12 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_13 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_14 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_15 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKINV_X2.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:47 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT CLKINV_X2 I ZN VDD VNW VPW VSS 
*.PININFO I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_i_0_0 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_1 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_1_0 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKINV_X20.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:53 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT CLKINV_X20 I ZN VDD VNW VPW VSS 
*.PININFO I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_i_0_0 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_1 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_2 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_3 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_4 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_5 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_6 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_7 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_8 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_9 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_10 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_11 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_12 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_13 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_14 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_15 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_16 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_17 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_18 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_19 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_1_0 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_4 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_5 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_6 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_7 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_8 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_9 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_10 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_11 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_12 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_13 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_14 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_15 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_16 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_17 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_18 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_19 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKINV_X3.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:48 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT CLKINV_X3 I ZN VDD VNW VPW VSS 
*.PININFO I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_i_0_0 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_1 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_2 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_1_0 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKINV_X4.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:48:46 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT CLKINV_X4 I ZN VDD VNW VPW VSS 
*.PININFO I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_i_0_0 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_1 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_2 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_3 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_1_0 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   CLKINV_X8.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:48:48 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT CLKINV_X8 I ZN VDD VNW VPW VSS 
*.PININFO I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_i_0_0_x8_0 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_0_x8_1 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_0_x8_2 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_0_x8_3 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_0_x8_4 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_0_x8_5 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_0_x8_6 ZN I VSS VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_0_0_x8_7 VSS I ZN VPW nmos_5p0 W=0.730000U L=0.600000U
M_i_1_0_x8_0 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0_x8_1 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0_x8_2 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0_x8_3 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0_x8_4 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0_x8_5 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0_x8_6 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0_x8_7 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFNQ_X1.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:47:22 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFNQ_X1 D CLKN Q VDD VNW VPW VSS 
*.PININFO D:I CLKN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn9 ncki CLKN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn16 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 VSS D net2 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn11 net2 cki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn0 net5 ncki net11 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 VSS net10 net11 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 net10 net5 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn2 net0 ncki net10 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn3 net7 cki net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 VSS net1 net7 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn5 net1 net0 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn6 Q net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp9 ncki CLKN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp16 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp10 VDD D net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp11 net5 ncki net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp0 net4 cki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp1 VDD net10 net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp15 net10 net5 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net0 cki net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net7 ncki net0 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 VDD net1 net7 VNW pmos_5p0 W=1.100000U L=0.500000U
M_tp3 net1 net0 VDD VNW pmos_5p0 W=1.100000U L=0.500000U
M_tp4 Q net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFNQ_X2.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:47:21 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFNQ_X2 D CLKN Q VDD VNW VPW VSS 
*.PININFO D:I CLKN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn9 ncki CLKN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn16 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 VSS D net2 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn11 net2 cki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn0 net5 ncki net11 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 VSS net10 net11 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 net10 net5 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn2 net0 ncki net10 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn3 net7 cki net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 VSS net1 net7 VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn5 net1 net0 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn6_7 Q net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn6 Q net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp9 ncki CLKN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp16 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp10 VDD D net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp11 net5 ncki net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp0 net4 cki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp1 VDD net10 net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp15 net10 net5 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net0 cki net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net7 ncki net0 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 VDD net1 net7 VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp3 net1 net0 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4_13 Q net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4 Q net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFNQ_X4.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs007             *
* at 11:47:18 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFNQ_X4 D CLKN Q VDD VNW VPW VSS 
*.PININFO D:I CLKN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn9 ncki CLKN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn16 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 VSS D net2 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn11 net2 cki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn0 net5 ncki net11 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 VSS net10 net11 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 net10 net5 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn2 net0 ncki net10 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn3 net7 cki net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 VSS net1 net7 VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn5 net1 net0 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn6_7 Q net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn6 Q net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn6_7_61 Q net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn6_49 Q net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp9 ncki CLKN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp16 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp10 VDD D net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp11 net5 ncki net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp0 net4 cki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp1 VDD net10 net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp15 net10 net5 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net0 cki net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net7 ncki net0 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 VDD net1 net7 VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp3 net1 net0 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4_13 Q net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4 Q net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4_13_64 Q net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4_55 Q net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFNRNQ_X1.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs007             *
* at 11:47:17 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFNRNQ_X1 D RN CLKN Q VDD VNW VPW VSS 
*.PININFO D:I RN:I CLKN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn13 ncki CLKN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn11 net6 D VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn15 net6 cki net1 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn14 net1 ncki net15 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn8 net12 net2 net15 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn9 VSS RN net12 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn18 VSS net1 net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn0 net8 ncki net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn1 net11 cki net8 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn12 net11 net4 VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn5 net0 RN VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn4 net4 net8 net0 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn3 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp11 ncki CLKN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp9 VDD D net6 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp15 net1 ncki net6 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net9 cki net1 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 VDD net2 net9 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net9 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 VDD net1 net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 net2 cki net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net8 ncki net11 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net11 net4 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net4 RN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp4 VDD net8 net4 VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp1 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFNRNQ_X2.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:47:16 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFNRNQ_X2 D RN CLKN Q VDD VNW VPW VSS 
*.PININFO D:I RN:I CLKN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn13 ncki CLKN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn11 net6 D VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn15 net6 cki net1 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn14 net1 ncki net15 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn8 net12 net2 net15 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn9 VSS RN net12 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn18 VSS net1 net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn0 net8 ncki net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn1 net11 cki net8 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn12 net11 net4 VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn5 net0 RN VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn4 net4 net8 net0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3_42 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp11 ncki CLKN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp9 VDD D net6 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp15 net1 ncki net6 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net9 cki net1 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 VDD net2 net9 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net9 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 VDD net1 net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 net2 cki net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net8 ncki net11 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net11 net4 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net4 RN VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4 VDD net8 net4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1_40 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFNRNQ_X4.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:47:19 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFNRNQ_X4 D RN CLKN Q VDD VNW VPW VSS 
*.PININFO D:I RN:I CLKN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn13 ncki CLKN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn11 net6 D VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn15 net6 cki net1 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn14 net1 ncki net15 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn8 net12 net2 net15 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn9 VSS RN net12 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn18 VSS net1 net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn0 net8 ncki net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn1 net11 cki net8 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn12 net11 net4 VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn5 net0 RN VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn4 net4 net8 net0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3_42 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3_42_63 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3_69 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp11 ncki CLKN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp9 VDD D net6 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp15 net1 ncki net6 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net9 cki net1 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 VDD net2 net9 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net9 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 VDD net1 net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 net2 cki net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net8 ncki net11 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net11 net4 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net4 RN VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4 VDD net8 net4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1_40 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1_40_64 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1_66 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFNRSNQ_X1.                                                     *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs010             *
* at 11:47:15 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFNRSNQ_X1 D RN SETN CLKN Q VDD VNW VPW VSS 
*.PININFO D:I RN:I SETN:I CLKN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn2 ncki CLKN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn1 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn0 net14 D VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn8 net14 cki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 net3 ncki net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net15 net4 net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn7 VSS RN net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn3 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net5 ncki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net7 cki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 net1 SETN net7 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn16 VSS net6 net1 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn18 net2 RN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn17 net6 net5 net2 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn19 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp2 ncki CLKN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp1 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp0 VDD D net14 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net3 ncki net14 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net13 cki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net13 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 VDD net3 net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp20 net4 cki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp19 net5 ncki net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 net7 SETN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp14 net7 net6 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp16 net6 RN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp15 VDD net5 net6 VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp17 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFNRSNQ_X2.                                                     *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs016             *
* at 11:47:16 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFNRSNQ_X2 D RN SETN CLKN Q VDD VNW VPW VSS 
*.PININFO D:I RN:I SETN:I CLKN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn2 ncki CLKN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn1 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn0 net14 D VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn8 net14 cki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 net3 ncki net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net15 net4 net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn7 VSS RN net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn3 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net5 ncki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net7 cki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 net1 SETN net7 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn16 VSS net6 net1 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn18 net2 RN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn17 net6 net5 net2 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn19_16 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn19 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp2 ncki CLKN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp1 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp0 VDD D net14 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net3 ncki net14 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net13 cki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net13 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 VDD net3 net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp20 net4 cki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp19 net5 ncki net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 net7 SETN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp14 net7 net6 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp16 net6 RN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp15 VDD net5 net6 VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp17_9 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp17 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFNRSNQ_X4.                                                     *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:47:16 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFNRSNQ_X4 D RN SETN CLKN Q VDD VNW VPW VSS 
*.PININFO D:I RN:I SETN:I CLKN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn2 ncki CLKN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn1 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn0 net14 D VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn8 net14 cki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 net3 ncki net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net15 net4 net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn7 VSS RN net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn3 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net5 ncki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net7 cki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 net1 SETN net7 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn16 VSS net6 net1 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn18 net2 RN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn17 net6 net5 net2 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn19_16 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn19 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn19_16_44 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn19_64 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp2 ncki CLKN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp1 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp0 VDD D net14 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net3 ncki net14 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net13 cki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net13 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 VDD net3 net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp20 net4 cki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp19 net5 ncki net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 net7 SETN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp14 net7 net6 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp16 net6 RN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp15 VDD net5 net6 VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp17_9 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp17 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp17_9_60 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp17_57 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFNSNQ_X1.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs027             *
* at 11:47:15 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFNSNQ_X1 D SETN CLKN Q VDD VNW VPW VSS 
*.PININFO D:I SETN:I CLKN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn0 ncki CLKN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn3 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 net13 D VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net13 cki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net3 ncki net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 VSS net4 net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn2 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net5 ncki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn12 net7 cki net5 VPW nmos_5p0 W=0.750000U L=0.600000U
M_tn14 net1 SETN net7 VPW nmos_5p0 W=0.750000U L=0.600000U
M_tn15 VSS net6 net1 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn18 net6 net5 VSS VPW nmos_5p0 W=0.750000U L=0.600000U
M_tn16 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp0 ncki CLKN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp4 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 VDD D net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 net3 ncki net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net10 cki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net4 net3 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 net5 cki net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp17 net7 ncki net5 VNW pmos_5p0 W=1.100000U L=0.500000U
M_tp12 net7 SETN VDD VNW pmos_5p0 W=1.100000U L=0.500000U
M_tp13 VDD net6 net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 net6 net5 VDD VNW pmos_5p0 W=1.100000U L=0.500000U
M_tp14 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFNSNQ_X2.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:47:14 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFNSNQ_X2 D SETN CLKN Q VDD VNW VPW VSS 
*.PININFO D:I SETN:I CLKN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn0 ncki CLKN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn3 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 net13 D VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net13 cki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net3 ncki net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 VSS net4 net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn2 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net5 ncki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn12 net7 cki net5 VPW nmos_5p0 W=0.750000U L=0.600000U
M_tn14 net1 SETN net7 VPW nmos_5p0 W=0.750000U L=0.600000U
M_tn15 VSS net6 net1 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn18 net6 net5 VSS VPW nmos_5p0 W=0.750000U L=0.600000U
M_tn16_30 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn16 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp0 ncki CLKN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp4 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 VDD D net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 net3 ncki net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net10 cki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net4 net3 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 net5 cki net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp17 net7 ncki net5 VNW pmos_5p0 W=1.100000U L=0.500000U
M_tp12 net7 SETN VDD VNW pmos_5p0 W=1.100000U L=0.500000U
M_tp13 VDD net6 net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 net6 net5 VDD VNW pmos_5p0 W=1.100000U L=0.500000U
M_tp14_24 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp14 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFNSNQ_X4.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:47:16 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFNSNQ_X4 D SETN CLKN Q VDD VNW VPW VSS 
*.PININFO D:I SETN:I CLKN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn0 ncki CLKN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn3 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 net13 D VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net13 cki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net3 ncki net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 VSS net4 net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn2 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net5 ncki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn12 net7 cki net5 VPW nmos_5p0 W=0.750000U L=0.600000U
M_tn14 net1 SETN net7 VPW nmos_5p0 W=0.750000U L=0.600000U
M_tn15 VSS net6 net1 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn18 net6 net5 VSS VPW nmos_5p0 W=0.750000U L=0.600000U
M_tn16_30 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn16 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn16_30_46 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn16_51 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp0 ncki CLKN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp4 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 VDD D net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 net3 ncki net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net10 cki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net4 net3 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 net5 cki net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp17 net7 ncki net5 VNW pmos_5p0 W=1.100000U L=0.500000U
M_tp12 net7 SETN VDD VNW pmos_5p0 W=1.100000U L=0.500000U
M_tp13 VDD net6 net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 net6 net5 VDD VNW pmos_5p0 W=1.100000U L=0.500000U
M_tp14_24 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp14 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp14_24_63 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp14_44 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFQ_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:47:09 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFQ_X1 D CLK Q VDD VNW VPW VSS 
*.PININFO D:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn3 VSS CLK ncki VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn4 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn5 net5 ncki VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn8 net4 D net5 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn6 net6 cki net4 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn7 VSS net0 net6 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn0 net0 net4 VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn9 net2 cki net0 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn11 net1 ncki net2 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn12 VSS net3 net1 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn10 net3 net2 VSS VPW nmos_5p0 W=0.750000U L=0.600000U
M_tn1 Q net3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp3 VDD CLK ncki VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp4 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp12 net7 cki VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp11 net4 D net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net8 ncki net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net0 net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp0 net0 net4 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net2 ncki net0 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 net1x cki net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 VDD net3 net1x VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp8 net3 net2 VDD VNW pmos_5p0 W=1.100000U L=0.500000U
M_tp1 Q net3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFQ_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:47:07 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFQ_X2 D CLK Q VDD VNW VPW VSS 
*.PININFO D:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn3 VSS CLK ncki VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn4 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn5 net5 ncki VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn8 net4 D net5 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn6 net6 cki net4 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn7 VSS net0 net6 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn0 net0 net4 VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn9 net2 cki net0 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn11 net1 ncki net2 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn12 VSS net3 net1 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn10 net3 net2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn1 Q net3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn1_18 Q net3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp3 VDD CLK ncki VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp4 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp12 net7 cki VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp11 net4 D net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net8 ncki net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net0 net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp0 net0 net4 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net2 ncki net0 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 net1x cki net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 VDD net3 net1x VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp8 net3 net2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1 Q net3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1_16 Q net3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFQ_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:47:08 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFQ_X4 D CLK Q VDD VNW VPW VSS 
*.PININFO D:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn3 VSS CLK ncki VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn4 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn5 net5 ncki VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn8 net4 D net5 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn6 net6 cki net4 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn7 VSS net0 net6 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn0 net0 net4 VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn9 net2 cki net0 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn11 net1 ncki net2 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn12 VSS net3 net1 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn10 net3 net2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn10_6 net3 net2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn1_39 Q net3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn1_18_47 Q net3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn1 Q net3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn1_18 Q net3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp3 VDD CLK ncki VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp4 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp12 net7 cki VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp11 net4 D net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net8 ncki net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net0 net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp0 net0 net4 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net2 ncki net0 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 net1x cki net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 VDD net3 net1x VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp8 net3 net2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp8_10 net3 net2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1_58 Q net3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1_16_34 Q net3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1 Q net3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1_16 Q net3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFRNQ_X1.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:47:09 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFRNQ_X1 D RN CLK Q VDD VNW VPW VSS 
*.PININFO D:I RN:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn10 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn13 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn11 net10 D VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn15 net10 ncki net1 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn14 net1 cki net15 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn8 net12 net2 net15 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn9 VSS RN net12 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn18 VSS net1 net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn0 net8 cki net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn1 net11 ncki net8 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn12 net11 net4 VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn5 net0 RN VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn4 net4 net8 net0 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn3 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp8 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp11 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp9 VDD D net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp15 net1 cki net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net9 ncki net1 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 VDD net2 net9 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net9 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 VDD net1 net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 net2 ncki net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net8 cki net11 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net11 net4 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net4 RN VDD VNW pmos_5p0 W=0.980000U L=0.500000U
M_tp4 VDD net8 net4 VNW pmos_5p0 W=0.980000U L=0.500000U
M_tp1 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFRNQ_X2.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs008             *
* at 11:47:07 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFRNQ_X2 D RN CLK Q VDD VNW VPW VSS 
*.PININFO D:I RN:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn10 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn13 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn11 net10 D VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn15 net10 ncki net1 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn14 net1 cki net15 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn8 net12 net2 net15 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn9 VSS RN net12 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn18 VSS net1 net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn0 net8 cki net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn1 net11 ncki net8 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn12 net11 net4 VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn5 net0 RN VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn4 net4 net8 net0 VPW nmos_5p0 W=1.180000U L=0.600000U
M_tn3_15 Q net4 VSS VPW nmos_5p0 W=1.250000U L=0.600000U
M_tn3 Q net4 VSS VPW nmos_5p0 W=1.250000U L=0.600000U
M_tp8 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp11 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp9 VDD D net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp15 net1 cki net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net9 ncki net1 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 VDD net2 net9 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net9 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 VDD net1 net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 net2 ncki net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net8 cki net11 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net11 net4 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net4 RN VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4 VDD net8 net4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1_13 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFRNQ_X4.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:47:09 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFRNQ_X4 D RN CLK Q VDD VNW VPW VSS 
*.PININFO D:I RN:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn10 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn13 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn11 net10 D VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 net10 ncki net1 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net1 cki net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn8 net12 net2 net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn9 VSS RN net12 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn18 VSS net1 net2 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn0 net8 cki net2 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 net11 ncki net8 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn12 net11 net4 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 net0 RN VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net4 net8 net0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3_15 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3_15_13 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3_10 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp8 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp11 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp9 VDD D net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp15 net1 cki net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net9 ncki net1 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 VDD net2 net9 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net9 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 VDD net1 net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 net2 ncki net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net8 cki net11 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net11 net4 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net4 RN VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4 VDD net8 net4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1_13 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1_13_25 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1_30 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFRSNQ_X1.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:47:11 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFRSNQ_X1 D RN SETN CLK Q VDD VNW VPW VSS 
*.PININFO D:I RN:I SETN:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn1 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn2 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn0 net14 D VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn8 net14 ncki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 net3 cki net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net15 net4 net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn7 VSS RN net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn3 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net5 cki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net7 ncki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 net1 SETN net7 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn16 VSS net6 net1 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn18 net2 RN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn17 net6 net5 net2 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn19 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp1 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp2 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp0 VDD D net14 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net3 cki net14 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net13 ncki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net13 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 VDD net3 net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp20 net4 ncki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp19 net5 cki net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 net7 SETN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp14 net7 net6 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp16 net6 RN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp15 VDD net5 net6 VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp17 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFRSNQ_X2.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs008             *
* at 11:47:06 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFRSNQ_X2 D RN SETN CLK Q VDD VNW VPW VSS 
*.PININFO D:I RN:I SETN:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn1 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn2 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn0 net14 D VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn8 net14 ncki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 net3 cki net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net15 net4 net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn7 VSS RN net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn3 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net5 cki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net7 ncki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 net1 SETN net7 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn16 VSS net6 net1 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn18 net2 RN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn17 net6 net5 net2 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn19_39 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn19 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp1 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp2 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp0 VDD D net14 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net3 cki net14 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net13 ncki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net13 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 VDD net3 net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp20 net4 ncki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp19 net5 cki net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 net7 SETN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp14 net7 net6 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp16 net6 RN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp15 VDD net5 net6 VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp17_33 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp17 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFRSNQ_X4.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs021             *
* at 11:47:09 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFRSNQ_X4 D RN SETN CLK Q VDD VNW VPW VSS 
*.PININFO D:I RN:I SETN:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn1 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn2 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn0 net14 D VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn8 net14 ncki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 net3 cki net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net15 net4 net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn7 VSS RN net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn3 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net5 cki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net7 ncki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 net1 SETN net7 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn16 VSS net6 net1 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn18 net2 RN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn17 net6 net5 net2 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn19_39 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn19 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn19_39_20 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn19_24 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp1 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp2 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp0 VDD D net14 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net3 cki net14 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net13 ncki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net13 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 VDD net3 net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp20 net4 ncki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp19 net5 cki net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 net7 SETN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp14 net7 net6 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp16 net6 RN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp15 VDD net5 net6 VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp17_33 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp17 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp17_33_0 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp17_16 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFSNQ_X1.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:47:07 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFSNQ_X1 D SETN CLK Q VDD VNW VPW VSS 
*.PININFO D:I SETN:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn3 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn0 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 net13 D VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net13 ncki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net3 cki net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 VSS net4 net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn2 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net5 cki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn12 net7 ncki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net1 SETN net7 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 VSS net6 net1 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn18 net6 net5 VSS VPW nmos_5p0 W=0.750000U L=0.600000U
M_tn16 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp4 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp0 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 VDD D net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 net3 cki net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net10 ncki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net4 net3 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 net5 ncki net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp17 net7 cki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net7 SETN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 VDD net6 net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 net6 net5 VDD VNW pmos_5p0 W=1.100000U L=0.500000U
M_tp14 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFSNQ_X2.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:47:08 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFSNQ_X2 D SETN CLK Q VDD VNW VPW VSS 
*.PININFO D:I SETN:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn3 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn0 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 net13 D VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net13 ncki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net3 cki net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 VSS net4 net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn2 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net5 cki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn12 net7 ncki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net1 SETN net7 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 VSS net6 net1 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn18 net6 net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn16 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn16_7 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp4 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp0 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 VDD D net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 net3 cki net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net10 ncki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net4 net3 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 net5 ncki net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp17 net7 cki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net7 SETN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 VDD net6 net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 net6 net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp14 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp14_2 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DFFSNQ_X4.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:47:08 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DFFSNQ_X4 D SETN CLK Q VDD VNW VPW VSS 
*.PININFO D:I SETN:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn3 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn0 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 net13 D VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net13 ncki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net3 cki net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 VSS net4 net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn2 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net5 cki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn12 net7 ncki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net1 SETN net7 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 VSS net6 net1 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn18 net6 net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn18_45 net6 net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn16 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn16_7 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn16_23 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn16_7_36 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp4 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp0 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 VDD D net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 net3 cki net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net10 ncki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net4 net3 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 net5 ncki net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp17 net7 cki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net7 SETN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 VDD net6 net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 net6 net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp16_52 net6 net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp14 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp14_2 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp14_19 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp14_2_27 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DLYA_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:44 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DLYA_X1 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 VSS Z_neg net_2 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_6 net_3 net_2 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_18 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1 VDD Z_neg net_2 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_29 net_3 net_2 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_3_0_0 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DLYA_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:45 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DLYA_X2 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 VSS Z_neg net_2 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_6 net_3 net_2 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_18 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0_18_1 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1 VDD Z_neg net_2 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_29 net_3 net_2 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_3_0_0 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0_0_14 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DLYA_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:44 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DLYA_X4 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 VSS Z_neg net_2 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_6 net_3 net_2 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_18 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0_18_1 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0_18_2 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0_18_1_15 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1 VDD Z_neg net_2 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_29 net_3 net_2 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_3_0_0 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0_0_14 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0_0_34 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0_0_14_19 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DLYB_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:43 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DLYB_X1 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 net_2 Z_neg net_1 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3 net_1 Z_neg VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_21 net_3 net_2 net_6 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_6 net_6 net_2 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_18 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0 net_0 Z_neg VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1 net_2 Z_neg net_0 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_29 net_5 net_2 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_39 net_3 net_2 net_5 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_3_0_0 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DLYB_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:45 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DLYB_X2 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 net_2 Z_neg net_1 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3 net_1 Z_neg VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_21 net_3 net_2 net_6 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_6 net_6 net_2 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_18 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0_18_1 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0 net_0 Z_neg VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1 net_2 Z_neg net_0 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_29 net_5 net_2 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_39 net_3 net_2 net_5 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_3_0_0 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0_0_14 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DLYB_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:48:43 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DLYB_X4 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 net_2 Z_neg net_1 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3 net_1 Z_neg VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_21 net_3 net_2 net_6 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_6 net_6 net_2 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_18 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0_18_1 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0_18_2 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0_18_1_15 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0 net_0 Z_neg VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1 net_2 Z_neg net_0 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_29 net_5 net_2 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_39 net_3 net_2 net_5 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_3_0_0 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0_0_14 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0_0_34 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0_0_14_19 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DLYC_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:45 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DLYC_X1 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 net_7 Z_neg net_1 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3 net_1 Z_neg VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_26 net_9 net_7 net_13 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_30 net_13 net_7 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_0 net_8 net_9 net_11 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_4 net_11 net_9 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_21 net_3 net_8 net_6 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_6 net_6 net_8 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_18 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0 net_0 Z_neg VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1 net_7 Z_neg net_0 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_35 net_12 net_7 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_47 net_9 net_7 net_12 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_9 net_10 net_9 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_22 net_8 net_9 net_10 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_29 net_5 net_8 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_39 net_3 net_8 net_5 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_3_0_0 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DLYC_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs016             *
* at 11:48:42 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DLYC_X2 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 net_7 Z_neg net_1 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3 net_1 Z_neg VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_26 net_9 net_7 net_13 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_30 net_13 net_7 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_0 net_8 net_9 net_11 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_4 net_11 net_9 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_21 net_3 net_8 net_6 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_6 net_6 net_8 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_18 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0_18_2 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0 net_0 Z_neg VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1 net_7 Z_neg net_0 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_35 net_12 net_7 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_47 net_9 net_7 net_12 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_9 net_10 net_9 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_22 net_8 net_9 net_10 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_29 net_5 net_8 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_39 net_3 net_8 net_5 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_3_0_0 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0_0_16 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DLYC_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:48:43 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DLYC_X4 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 net_7 Z_neg net_1 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3 net_1 Z_neg VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_26 net_9 net_7 net_13 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_30 net_13 net_7 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_0 net_8 net_9 net_11 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_4 net_11 net_9 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_21 net_3 net_8 net_6 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_6 net_6 net_8 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_18 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0_18_2 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0_18_1 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0_18_2_36 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0 net_0 Z_neg VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1 net_7 Z_neg net_0 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_35 net_12 net_7 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_47 net_9 net_7 net_12 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_9 net_10 net_9 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_22 net_8 net_9 net_10 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_29 net_5 net_8 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_39 net_3 net_8 net_5 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_3_0_0 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0_0_16 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0_0_32 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0_0_16_16 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DLYD_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs027             *
* at 11:48:42 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DLYD_X1 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 net_7 Z_neg net_1 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3 net_1 Z_neg VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_26 net_9 net_7 net_13 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_30 net_13 net_7 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_0 net_15 net_9 net_11 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_4 net_11 net_9 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_26_13 net_16 net_15 net_18 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_30_34 net_18 net_15 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_10 net_14 net_16 net_19 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_4_49 net_19 net_16 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_21 net_3 net_14 net_6 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_6 net_6 net_14 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_18 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0 net_0 Z_neg VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1 net_7 Z_neg net_0 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_35 net_12 net_7 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_47 net_9 net_7 net_12 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_9 net_10 net_9 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_22 net_15 net_9 net_10 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_35_50 net_17 net_15 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_47_46 net_16 net_15 net_17 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_9_2 net_20 net_16 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_22_38 net_14 net_16 net_20 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_29 net_5 net_14 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_39 net_3 net_14 net_5 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_3_0_0 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DLYD_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:44 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DLYD_X2 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 net_7 Z_neg net_1 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3 net_1 Z_neg VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_26 net_9 net_7 net_13 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_30 net_13 net_7 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_0 net_15 net_9 net_11 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_4 net_11 net_9 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_26_13 net_16 net_15 net_18 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_30_34 net_18 net_15 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_10 net_14 net_16 net_19 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_4_49 net_19 net_16 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_21 net_3 net_14 net_6 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_6 net_6 net_14 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_18 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0_18_1 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0 net_0 Z_neg VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1 net_7 Z_neg net_0 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_35 net_12 net_7 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_47 net_9 net_7 net_12 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_9 net_10 net_9 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_22 net_15 net_9 net_10 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_35_50 net_17 net_15 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_47_46 net_16 net_15 net_17 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_9_2 net_20 net_16 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_22_38 net_14 net_16 net_20 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_29 net_5 net_14 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_39 net_3 net_14 net_5 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_3_0_0 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0_0_14 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   DLYD_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:48:44 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT DLYD_X4 I Z VDD VNW VPW VSS 
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 net_7 Z_neg net_1 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3 net_1 Z_neg VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_26 net_9 net_7 net_13 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_30 net_13 net_7 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_0 net_15 net_9 net_11 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_4 net_11 net_9 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_26_13 net_16 net_15 net_18 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_30_34 net_18 net_15 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_10 net_14 net_16 net_19 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_4_49 net_19 net_16 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_21 net_3 net_14 net_6 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_3_6 net_6 net_14 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2_0_18 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0_18_1 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0_18_2 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0_18_1_15 Z net_3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0 net_0 Z_neg VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1 net_7 Z_neg net_0 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_35 net_12 net_7 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_47 net_9 net_7 net_12 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_9 net_10 net_9 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_22 net_15 net_9 net_10 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_35_50 net_17 net_15 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_47_46 net_16 net_15 net_17 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_9_2 net_20 net_16 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_22_38 net_14 net_16 net_20 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_0_29 net_5 net_14 VDD VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_1_39 net_3 net_14 net_5 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_3_0_0 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0_0_14 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0_0_34 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0_0_14_19 Z net_3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FILLCAP_X16.                                                     *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:48:59 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT FILLCAP_X16 VDD VNW VPW VSS 
*.PININFO VDD:P VNW:P VPW:P VSS:G 
M_i_17 net_3 net_2 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_23 net_4 net_5 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_24 net_7 net_9 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_23_55 net_6 net_8 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_19 VDD net_3 net_2 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_7 VDD net_4 net_5 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_33 VDD net_7 net_9 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_7_23 VDD net_6 net_8 VNW pmos_5p0 W=1.830000U L=1.000000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FILLCAP_X32.                                                     *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:49:04 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT FILLCAP_X32 VDD VNW VPW VSS 
*.PININFO VDD:P VNW:P VPW:P VSS:G 
M_i_17 net_3 net_2 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_23 net_4 net_5 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_24 net_7 net_9 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_23_55 net_6 net_8 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_27 net_17 net_14 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_23_63 net_16 net_15 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_24_22 net_13 net_11 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_23_55_93 net_12 net_10 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_19 VDD net_3 net_2 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_7 VDD net_4 net_5 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_33 VDD net_7 net_9 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_7_23 VDD net_6 net_8 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_94 VDD net_17 net_14 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_7_87 VDD net_16 net_15 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_33_95 VDD net_13 net_11 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_7_23_23 VDD net_12 net_10 VNW pmos_5p0 W=1.830000U L=1.000000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FILLCAP_X4.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:49:00 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT FILLCAP_X4 VDD VNW VPW VSS 
*.PININFO VDD:P VNW:P VPW:P VSS:G 
M_i_17 net_1 net_0 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_19 VDD net_1 net_0 VNW pmos_5p0 W=1.830000U L=1.000000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FILLCAP_X64.                                                     *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:49:08 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT FILLCAP_X64 VDD VNW VPW VSS 
*.PININFO VDD:P VNW:P VPW:P VSS:G 
M_i_17 net_3 net_2 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_23 net_4 net_5 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_24 net_7 net_9 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_23_55 net_6 net_8 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_27 net_17 net_14 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_23_63 net_16 net_15 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_24_22 net_13 net_11 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_23_55_93 net_12 net_10 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_20 net_30 net_26 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_23_59 net_25 net_20 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_24_135 net_23 net_28 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_23_55_90 net_33 net_18 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_27_139 net_31 net_29 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_23_63_82 net_32 net_24 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_24_22_30 net_22 net_27 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_23_55_93_110 net_19 net_21 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_19 VDD net_3 net_2 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_7 VDD net_4 net_5 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_33 VDD net_7 net_9 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_7_23 VDD net_6 net_8 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_94 VDD net_17 net_14 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_7_87 VDD net_16 net_15 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_33_95 VDD net_13 net_11 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_7_23_23 VDD net_12 net_10 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_95 VDD net_30 net_26 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_7_188 VDD net_25 net_20 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_33_98 VDD net_23 net_28 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_7_23_16 VDD net_33 net_18 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_94_91 VDD net_31 net_29 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_7_87_65 VDD net_32 net_24 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_33_95_109 VDD net_22 net_27 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_7_23_23_99 VDD net_19 net_21 VNW pmos_5p0 W=1.830000U L=1.000000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FILLCAP_X8.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:49:00 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT FILLCAP_X8 VDD VNW VPW VSS 
*.PININFO VDD:P VNW:P VPW:P VSS:G 
M_i_17 net_3 net_2 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_23 net_4 net_5 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_19 VDD net_3 net_2 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_7 VDD net_4 net_5 VNW pmos_5p0 W=1.830000U L=1.000000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FILLTIE.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:49:01 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT FILLTIE VDD VSS 
*.PININFO VDD:P VSS:G 
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   HOLD.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs016             *
* at 11:49:00 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT HOLD Z VDD VNW VPW VSS 
*.PININFO Z:B VDD:P VNW:P VPW:P VSS:G 
M_u7 VDD Z net8 VNW pmos_5p0 W=1.830000U L=0.500000U
M_u3 VSS Z net8 VPW nmos_5p0 W=1.320000U L=0.600000U
M_MU12 Z net8 VDD VNW pmos_5p0 W=0.360000U L=2.00000U
M_MU11 Z net8 VSS VPW nmos_5p0 W=0.360000U L=2.00000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   ICGTN_X1.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:47:01 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT ICGTN_X1 CLKN E TE Q VDD VNW VPW VSS 
*.PININFO CLKN:I E:I TE:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_MU19 VSS TE net50 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU20 net50 E VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI82 net53 NCP net50 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI91 net038 CP net53 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI92 VSS QD net038 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU82_M_u2 NCP CP VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI95_M_u2 VSS net53 QD VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI89_M_u2 net36 QD VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU81_M_u2 VSS CLKN CP VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI1_M_u3 d3 net36 VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI1_M_u4 VSS CLKN d3 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU75_M_u2 Q d3 VSS VPW nmos_5p0 W=1.000000U L=0.600000U
M_MI81 net58 TE VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU17 net61 E net58 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU16 net53 CP net61 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI90 net067 NCP net53 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI88 VDD QD net067 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU82_M_u3 NCP CP VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI95_M_u3 VDD net53 QD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI89_M_u3 net36 QD VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU81_M_u3 VDD CLKN CP VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI1_M_u1 XI1-net8 net36 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI1_M_u2 d3 CLKN XI1-net8 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU75_M_u3 Q d3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   ICGTN_X2.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:46:59 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT ICGTN_X2 CLKN E TE Q VDD VNW VPW VSS 
*.PININFO CLKN:I E:I TE:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_MU19 VSS TE net50 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU20 net50 E VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI82 net53 NCP net50 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI91 net038 CP net53 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI92 VSS QD net038 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU82_M_u2 NCP CP VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI95_M_u2 VSS net53 QD VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI89_M_u2 net36 QD VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU81_M_u2 VSS CLKN CP VPW nmos_5p0 W=0.800000U L=0.600000U
M_MI1_M_u3 d3 net36 VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_MI1_M_u4 VSS CLKN d3 VPW nmos_5p0 W=0.800000U L=0.600000U
M_MU75_M_u2 Q d3 VSS VPW nmos_5p0 W=1.000000U L=0.600000U
M_MU75_M_u2_19 Q d3 VSS VPW nmos_5p0 W=1.000000U L=0.600000U
M_MI81 net58 TE VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU17 net61 E net58 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU16 net53 CP net61 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI90 net067 NCP net53 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI88 VDD QD net067 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU82_M_u3 NCP CP VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI95_M_u3 VDD net53 QD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI89_M_u3 net36 QD VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU81_M_u3 VDD CLKN CP VNW pmos_5p0 W=1.680000U L=0.500000U
M_MI1_M_u1 XI1-net8 net36 VDD VNW pmos_5p0 W=1.680000U L=0.500000U
M_MI1_M_u2 d3 CLKN XI1-net8 VNW pmos_5p0 W=1.680000U L=0.500000U
M_MU75_M_u3 Q d3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_MU75_M_u3_1 Q d3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   ICGTN_X4.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:46:43 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT ICGTN_X4 CLKN E TE Q VDD VNW VPW VSS 
*.PININFO CLKN:I E:I TE:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_MU19 VSS TE net50 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU20 net50 E VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI82 net53 NCP net50 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI91 net038 CP net53 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI92 VSS QD net038 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU82_M_u2 NCP CP VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI95_M_u2 VSS net53 QD VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI89_M_u2 net36 QD VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU81_M_u2 VSS CLKN CP VPW nmos_5p0 W=0.800000U L=0.600000U
M_MI1_M_u3 d3 net36 VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_MI1_M_u4 VSS CLKN d3 VPW nmos_5p0 W=0.800000U L=0.600000U
M_MU75_M_u2 Q d3 VSS VPW nmos_5p0 W=1.000000U L=0.600000U
M_MU75_M_u2_19 Q d3 VSS VPW nmos_5p0 W=1.000000U L=0.600000U
M_MU75_M_u2_33 Q d3 VSS VPW nmos_5p0 W=1.000000U L=0.600000U
M_MU75_M_u2_19_5 Q d3 VSS VPW nmos_5p0 W=1.000000U L=0.600000U
M_MI81 net58 TE VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU17 net61 E net58 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU16 net53 CP net61 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI90 net067 NCP net53 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI88 VDD QD net067 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU82_M_u3 NCP CP VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI95_M_u3 VDD net53 QD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI89_M_u3 net36 QD VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU81_M_u3 VDD CLKN CP VNW pmos_5p0 W=1.680000U L=0.500000U
M_MI1_M_u1 XI1-net8 net36 VDD VNW pmos_5p0 W=1.680000U L=0.500000U
M_MI1_M_u2 d3 CLKN XI1-net8 VNW pmos_5p0 W=1.680000U L=0.500000U
M_MU75_M_u3 Q d3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_MU75_M_u3_1 Q d3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_MU75_M_u3_2 Q d3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_MU75_M_u3_1_35 Q d3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   ICGTP_X1.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:46:41 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT ICGTP_X1 CLK E TE Q VDD VNW VPW VSS 
*.PININFO CLK:I E:I TE:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_MU19 net50 TE VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU20 VSS E net50 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI82 net50 NCK net53 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI91 net53 CK net033 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI92 net033 QD VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI80_M_u2 VSS net53 QD VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU82_M_u2 VSS NCK CK VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU81_M_u2 NCK CLK VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI85_M_u3 XI85-net6 CLK d3 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI85_M_u4 VSS QD XI85-net6 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU75_M_u2 Q d3 VSS VPW nmos_5p0 W=1.000000U L=0.600000U
M_MI81 VDD TE net58 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU17 net58 E net61 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU16 net61 CK net53 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI90 net53 NCK net062 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI88 net062 QD VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI80_M_u3 VDD net53 QD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU82_M_u3 CK NCK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU81_M_u3 VDD CLK NCK VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI85_M_u1 d3 CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI85_M_u2 VDD QD d3 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU75_M_u3 Q d3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   ICGTP_X2.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:46:42 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT ICGTP_X2 CLK E TE Q VDD VNW VPW VSS 
*.PININFO CLK:I E:I TE:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_MU19 net50 TE VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU20 VSS E net50 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI82 net50 NCK net53 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI91 net53 CK net033 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI92 net033 QD VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI80_M_u2 VSS net53 QD VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU82_M_u2 VSS NCK CK VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU81_M_u2 NCK CLK VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI85_M_u3 XI85-net6 CLK d3 VPW nmos_5p0 W=1.000000U L=0.600000U
M_MI85_M_u4 VSS QD XI85-net6 VPW nmos_5p0 W=1.000000U L=0.600000U
M_MU75_M_u2 Q d3 VSS VPW nmos_5p0 W=1.000000U L=0.600000U
M_MU75_M_u2_22 Q d3 VSS VPW nmos_5p0 W=1.000000U L=0.600000U
M_MI81 VDD TE net58 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU17 net58 E net61 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU16 net61 CK net53 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI90 net53 NCK net062 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI88 net062 QD VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI80_M_u3 VDD net53 QD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU82_M_u3 CK NCK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU81_M_u3 VDD CLK NCK VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI85_M_u1 d3 CLK VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_MI85_M_u2 VDD QD d3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_MU75_M_u3 Q d3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_MU75_M_u3_3 Q d3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   ICGTP_X4.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:46:42 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT ICGTP_X4 CLK E TE Q VDD VNW VPW VSS 
*.PININFO CLK:I E:I TE:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_MU19 net50 TE VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU20 VSS E net50 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI82 net50 NCK net53 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI91 net53 CK net033 VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI92 net033 QD VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI80_M_u2 VSS net53 QD VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU82_M_u2 VSS NCK CK VPW nmos_5p0 W=0.700000U L=0.600000U
M_MU81_M_u2 NCK CLK VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_MI85_M_u3 XI85-net6 CLK d3 VPW nmos_5p0 W=1.000000U L=0.600000U
M_MI85_M_u4 VSS QD XI85-net6 VPW nmos_5p0 W=1.000000U L=0.600000U
M_MU75_M_u2 Q d3 VSS VPW nmos_5p0 W=1.000000U L=0.600000U
M_MU75_M_u2_22 Q d3 VSS VPW nmos_5p0 W=1.000000U L=0.600000U
M_MU75_M_u2_41 Q d3 VSS VPW nmos_5p0 W=1.000000U L=0.600000U
M_MU75_M_u2_22_37 Q d3 VSS VPW nmos_5p0 W=1.000000U L=0.600000U
M_MI81 VDD TE net58 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU17 net58 E net61 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU16 net61 CK net53 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI90 net53 NCK net062 VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI88 net062 QD VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI80_M_u3 VDD net53 QD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU82_M_u3 CK NCK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MU81_M_u3 VDD CLK NCK VNW pmos_5p0 W=1.380000U L=0.500000U
M_MI85_M_u1 d3 CLK VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_MI85_M_u2 VDD QD d3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_MU75_M_u3 Q d3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_MU75_M_u3_3 Q d3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_MU75_M_u3_1 Q d3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_MU75_M_u3_3_28 Q d3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INVZ_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:48:32 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT INVZ_X1 EN I ZN VDD VNW VPW VSS 
*.PININFO EN:I I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_mn VSS EN NEN VPW nmos_5p0 W=0.590000U L=0.600000U
M_mn8 NI_N NEN VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_mn21 NI_P EN NI_N VPW nmos_5p0 W=0.590000U L=0.600000U
M_mn3 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17 VSS NI NI_N VPW nmos_5p0 W=0.590000U L=0.600000U
M_Mn_inv NI I VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_mp VDD EN NEN VNW pmos_5p0 W=0.990000U L=0.500000U
M_mp7 NI_P EN VDD VNW pmos_5p0 W=0.990000U L=0.500000U
M_mp22 NI_N NEN NI_P VNW pmos_5p0 W=0.990000U L=0.500000U
M_mp4 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14 VDD NI NI_P VNW pmos_5p0 W=0.990000U L=0.500000U
M_Mp_inv NI I VDD VNW pmos_5p0 W=0.990000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INVZ_X12.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs024             *
* at 11:48:41 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT INVZ_X12 EN I ZN VDD VNW VPW VSS 
*.PININFO EN:I I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_mn VSS EN NEN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn8 NI_N NEN VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn21 NI_P EN NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_Mn_inv1 VSS I NI VPW nmos_5p0 W=1.320000U L=0.600000U
M_Mn_inv2 NI I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_Mn_inv3 VSS I NI VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17 NI_N NI VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9 VSS NI NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_10 NI_N NI VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9_17 VSS NI NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_10_0 NI_N NI VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9_17_30 VSS NI NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_89 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_34 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49_80 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25_35 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_99 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_33 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49_88 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25_34 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mp VDD EN NEN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp7 NI_P EN VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp22 NI_N NEN NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_Mp_inv1 VDD I NI VNW pmos_5p0 W=1.800000U L=0.500000U
M_Mp_inv2 NI I VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_Mp_inv3 VDD I NI VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14 NI_P NI VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10 VDD NI NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_11 NI_P NI VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10_8 VDD NI NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_11_21 NI_P NI VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10_8_17 VDD NI NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_57 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_96 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56_105 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57_69 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_58 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_106 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56_111 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57_75 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INVZ_X16.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:48:46 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT INVZ_X16 EN I ZN VDD VNW VPW VSS 
*.PININFO EN:I I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_mn VSS EN NEN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn8 NI_N NEN VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn21 NI_P EN NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_Mn_inv1 NI I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_Mn_inv2 VSS I NI VPW nmos_5p0 W=1.320000U L=0.600000U
M_Mn_inv3 NI I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_Mn_inv4 VSS I NI VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17 NI_N NI VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9 VSS NI NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_10 NI_N NI VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9_17 VSS NI NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_34 NI_N NI VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9_41 VSS NI NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_10_30 NI_N NI VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9_17_61 VSS NI NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_118 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_65 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49_181 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25_137 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_99_125 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_33_198 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49_88_82 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25_34_75 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_99 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_33 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49_88 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25_34 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mp VDD EN NEN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp7 NI_P EN VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp22 NI_N NEN NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_Mp_inv1 NI I VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_Mp_inv2 VDD I NI VNW pmos_5p0 W=1.800000U L=0.500000U
M_Mp_inv3 NI I VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_Mp_inv4 VDD I NI VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14 NI_P NI VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10 VDD NI NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_11 NI_P NI VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10_8 VDD NI NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_7 NI_P NI VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10_32 VDD NI NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_11_55 NI_P NI VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10_8_20 VDD NI NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_153 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_126 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56_133 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57_97 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_58_95 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_106_111 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56_111_134 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57_75_85 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_58 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_106 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56_111 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57_75 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INVZ_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs007             *
* at 11:48:30 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT INVZ_X2 EN I ZN VDD VNW VPW VSS 
*.PININFO EN:I I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_XX27 VSS EN NEN VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX44 NI_N NEN VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX36 NI_P EN NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX43 VSS NI NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX22 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX22_4 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_Mn_inv NI I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX28 VDD EN NEN VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX45 NI_P EN VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX39 NI_N NEN NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX46 VDD NI NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX21 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_XX21_5 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_Mp_inv NI I VDD VNW pmos_5p0 W=1.800000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INVZ_X3.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:48:31 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT INVZ_X3 EN I ZN VDD VNW VPW VSS 
*.PININFO EN:I I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_mn VSS EN NEN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn8 NI_N NEN VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn21 NI_P EN NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_Mn_inv VSS I NI VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17 NI_N NI VSS VPW nmos_5p0 W=0.885000U L=0.600000U
M_mn17_1 VSS NI NI_N VPW nmos_5p0 W=0.885000U L=0.600000U
M_mn3 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_2 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mp VDD EN NEN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp7 NI_P EN VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp22 NI_N NEN NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_Mp_inv VDD I NI VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14 NI_P NI VDD VNW pmos_5p0 W=1.485000U L=0.500000U
M_mp14_1 VDD NI NI_P VNW pmos_5p0 W=1.485000U L=0.500000U
M_mp4 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_1 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_2 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INVZ_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:48:30 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT INVZ_X4 EN I ZN VDD VNW VPW VSS 
*.PININFO EN:I I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_mn VSS EN NEN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn8 NI_N NEN VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn21 NI_P EN NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_Mn_inv VSS I NI VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17 NI_N NI VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9 VSS NI NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mp VDD EN NEN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp7 NI_P EN VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp22 NI_N NEN NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_Mp_inv VDD I NI VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14 NI_P NI VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10 VDD NI NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INVZ_X8.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:48:33 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT INVZ_X8 EN I ZN VDD VNW VPW VSS 
*.PININFO EN:I I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_mn VSS EN NEN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn8 NI_N NEN VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn21 NI_P EN NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_Mn_inv1 NI I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_Mn_inv2 VSS I NI VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17 NI_N NI VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9 VSS NI NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_10 NI_N NI VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn17_9_17 VSS NI NI_N VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_99 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_33 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_49_88 ZN NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_mn3_1_25_34 VSS NI_N ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_mp VDD EN NEN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp7 NI_P EN VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp22 NI_N NEN NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_Mp_inv1 NI I VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_Mp_inv2 VDD I NI VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14 NI_P NI VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10 VDD NI NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_11 NI_P NI VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp14_10_8 VDD NI NI_P VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_58 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_106 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_56_111 ZN NI_P VDD VNW pmos_5p0 W=1.800000U L=0.500000U
M_mp4_12_57_75 VDD NI_P ZN VNW pmos_5p0 W=1.800000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INV_X1.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:48:36 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT INV_X1 I ZN VDD VNW VPW VSS 
*.PININFO I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_i_0 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INV_X12.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:48:38 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT INV_X12 I ZN VDD VNW VPW VSS 
*.PININFO I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_i_0_0 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_4 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_5 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_6 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_7 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_8 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_9 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_10 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_11 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_4 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_5 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_6 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_7 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_8 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_9 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_10 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_11 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INV_X16.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:41 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT INV_X16 I ZN VDD VNW VPW VSS 
*.PININFO I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_i_0_0 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_4 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_5 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_6 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_7 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_8 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_9 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_10 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_11 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_12 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_13 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_14 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_15 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_4 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_5 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_6 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_7 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_8 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_9 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_10 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_11 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_12 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_13 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_14 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_15 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INV_X2.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs024             *
* at 11:48:37 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT INV_X2 I ZN VDD VNW VPW VSS 
*.PININFO I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_i_0_0 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INV_X20.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:44 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT INV_X20 I ZN VDD VNW VPW VSS 
*.PININFO I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_i_0_0 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_4 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_5 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_6 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_7 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_8 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_9 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_10 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_11 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_12 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_13 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_14 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_15 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_16 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_17 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_18 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_19 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_4 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_5 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_6 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_7 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_8 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_9 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_10 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_11 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_12 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_13 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_14 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_15 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_16 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_17 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_18 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_19 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INV_X3.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:36 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT INV_X3 I ZN VDD VNW VPW VSS 
*.PININFO I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_i_0_0 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INV_X4.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs021             *
* at 11:48:36 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT INV_X4 I ZN VDD VNW VPW VSS 
*.PININFO I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_i_0_0 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   INV_X8.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs007             *
* at 11:48:36 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT INV_X8 I ZN VDD VNW VPW VSS 
*.PININFO I:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!I
M_i_0_0_x8_0 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0_x8_1 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0_x8_2 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0_x8_3 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0_x8_4 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0_x8_5 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0_x8_6 ZN I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0_x8_7 VSS I ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0_x8_0 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0_x8_1 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0_x8_2 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0_x8_3 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0_x8_4 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0_x8_5 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0_x8_6 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0_x8_7 VDD I ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   LATQ_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:46:40 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT LATQ_X1 D E Q VDD VNW VPW VSS 
*.PININFO D:I E:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn0 VSS E net4 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn8 net7 net4 VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn4 VSS D net3 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn5 net5 net7 net3 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn1 net2 net4 net5 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn2 net2 net6 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn3 net6 net5 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn6 Q net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp0 VDD E net4 VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 net7 net4 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD D net1 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 net1 net4 net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 net5 net7 net0 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp1 net0 net6 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp3 net6 net5 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp6 Q net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   LATQ_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs021             *
* at 11:46:40 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT LATQ_X2 D E Q VDD VNW VPW VSS 
*.PININFO D:I E:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn0 VSS E net4 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn8 net7 net4 VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn4 VSS D net3 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn5 net5 net7 net3 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn1 net2 net4 net5 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn2 net2 net6 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn3 net6 net5 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn6_30 Q net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn6 Q net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp0 VDD E net4 VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 net7 net4 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD D net1 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 net1 net4 net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 net5 net7 net0 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp1 net0 net6 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp3 net6 net5 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp6_31 Q net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp6 Q net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   LATQ_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:46:39 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT LATQ_X4 D E Q VDD VNW VPW VSS 
*.PININFO D:I E:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn0 VSS E net4 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn8 net7 net4 VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn4 VSS D net3 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn5 net5 net7 net3 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn1 net2 net4 net5 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn2 net2 net6 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn3 net6 net5 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn3_94 net6 net5 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn6_30_66 Q net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn6_46 Q net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn6_30 Q net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn6 Q net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp0 VDD E net4 VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 net7 net4 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD D net1 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 net1 net4 net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 net5 net7 net0 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp1 net0 net6 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp3 net6 net5 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp3_85 net6 net5 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp6_31_68 Q net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp6_71 Q net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp6_31 Q net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp6 Q net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   LATRNQ_X1.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:46:38 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT LATRNQ_X1 D E RN Q VDD VNW VPW VSS 
*.PININFO D:I E:I RN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn3 net7 E VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 net1 RN VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn9 net2 D net1 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn8 net2 E net3 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn7 net3 net7 net4 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn5 net5 net0 net4 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn0 VSS RN net5 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn6 net0 net3 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn4 net6 net0 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn1 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp2 net7 E VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 VDD RN net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net8 D VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net3 net7 net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 net9 E net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net9 net0 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 net0 net3 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp7 net6 net0 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp0 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   LATRNQ_X2.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:46:38 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT LATRNQ_X2 D E RN Q VDD VNW VPW VSS 
*.PININFO D:I E:I RN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn3 net7 E VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 net1 RN VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn9 net2 D net1 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn8 net2 E net3 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn7 net3 net7 net4 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn5 net5 net0 net4 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn0 VSS RN net5 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn6 net0 net3 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn4 net6 net0 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn1 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn1_38 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp2 net7 E VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 VDD RN net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net8 D VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net3 net7 net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 net9 E net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net9 net0 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 net0 net3 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp7 net6 net0 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp0 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp0_27 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   LATRNQ_X4.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:46:40 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT LATRNQ_X4 D E RN Q VDD VNW VPW VSS 
*.PININFO D:I E:I RN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn3 net7 E VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 net1 RN VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn9 net2 D net1 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn8 net2 E net3 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn7 net3 net7 net4 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn5 net5 net0 net4 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn0 VSS RN net5 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn6 net0 net3 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn6_109 net0 net3 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn4 net6 net0 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn4_77 net6 net0 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn1 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn1_38 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn1_15 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn1_38_14 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp2 net7 E VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 VDD RN net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net8 D VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net3 net7 net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 net9 E net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net9 net0 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 net0 net3 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp9_110 net0 net3 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp7 net6 net0 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp7_78 net6 net0 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp0 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp0_27 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp0_24 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp0_27_20 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   LATRSNQ_X1.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:46:39 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT LATRSNQ_X1 D E RN SETN Q VDD VNW VPW VSS 
*.PININFO D:I E:I RN:I SETN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn3 net8 E VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn9 net2 RN VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn8 net3 D net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn7 net3 E net4 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn6 net4 net8 net5 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn5 net6 net1 net5 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn0 VSS RN net6 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn11 VSS net4 net0 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 net0 SETN net1 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn4 net7 net1 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn1 Q net7 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp2 net8 E VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 VDD RN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net9 D VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net4 net8 net9 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 net10 E net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net10 net1 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 VDD net4 net1 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 net1 SETN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp7 net7 net1 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp0 Q net7 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   LATRSNQ_X2.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:46:38 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT LATRSNQ_X2 D E RN SETN Q VDD VNW VPW VSS 
*.PININFO D:I E:I RN:I SETN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn3 net8 E VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn9 net2 RN VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn8 net3 D net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn7 net3 E net4 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn6 net4 net8 net5 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn5 net6 net1 net5 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn0 VSS RN net6 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn11 VSS net4 net0 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 net0 SETN net1 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn4 net7 net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn1 Q net7 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn1_19 Q net7 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp2 net8 E VDD VNW pmos_5p0 W=1.380000U L=0.600000U
M_tp8 VDD RN net4 VNW pmos_5p0 W=1.000000U L=0.600000U
M_tp6 net9 D VDD VNW pmos_5p0 W=1.000000U L=0.600000U
M_tp5 net4 net8 net9 VNW pmos_5p0 W=1.000000U L=0.600000U
M_tp4 net10 E net4 VNW pmos_5p0 W=1.000000U L=0.600000U
M_tp3 net10 net1 VDD VNW pmos_5p0 W=1.000000U L=0.600000U
M_tp10 VDD net4 net1 VNW pmos_5p0 W=1.000000U L=0.600000U
M_tp9 net1 SETN VDD VNW pmos_5p0 W=1.380000U L=0.600000U
M_tp7 net7 net1 VDD VNW pmos_5p0 W=1.830000U L=0.600000U
M_tp0 Q net7 VDD VNW pmos_5p0 W=1.830000U L=0.600000U
M_tp0_9 Q net7 VDD VNW pmos_5p0 W=1.830000U L=0.600000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   LATRSNQ_X4.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:46:40 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT LATRSNQ_X4 D E RN SETN Q VDD VNW VPW VSS 
*.PININFO D:I E:I RN:I SETN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn3 net8 E VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn9 net2 RN VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn8 net3 D net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn7 net3 E net4 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn6 net4 net8 net5 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn5 net6 net1 net5 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn0 VSS RN net6 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn11 VSS net4 net0 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 net0 SETN net1 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn4_44 net7 net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn4 net7 net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn1 Q net7 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn1_19 Q net7 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn1_18 Q net7 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn1_19_0 Q net7 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp2 net8 E VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 VDD RN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net9 D VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net4 net8 net9 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 net10 E net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net10 net1 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 VDD net4 net1 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 net1 SETN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp7_47 net7 net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp7 net7 net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp0 Q net7 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp0_9 Q net7 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp0_26 Q net7 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp0_9_34 Q net7 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   LATSNQ_X1.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:46:37 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT LATSNQ_X1 D E SETN Q VDD VNW VPW VSS 
*.PININFO D:I E:I SETN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn2 net6 E VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn7 VSS D net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn6 net3 E net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn5 net4 net6 net3 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn4 net4 net1 VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn9 VSS net3 net0 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn8 net0 SETN net1 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn3 net5 net1 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn0 Q net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp2 net6 E VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp6 VDD D net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net7 net6 net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 net3 E net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net8 net1 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 VDD net3 net1 VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 net1 SETN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp7 net5 net1 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp0 Q net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   LATSNQ_X2.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:46:37 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT LATSNQ_X2 D E SETN Q VDD VNW VPW VSS 
*.PININFO D:I E:I SETN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn2 net6 E VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn7 VSS D net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn6 net3 E net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn5 net4 net6 net3 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn4 net4 net1 VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn9 VSS net3 net0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn8 net0 SETN net1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3 net5 net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn0 Q net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn0_11 Q net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp2 net6 E VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp6 VDD D net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net7 net6 net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 net3 E net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net8 net1 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 VDD net3 net1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp8 net1 SETN VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp7 net5 net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp0 Q net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp0_8 Q net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   LATSNQ_X4.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:46:38 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT LATSNQ_X4 D E SETN Q VDD VNW VPW VSS 
*.PININFO D:I E:I SETN:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn2 net6 E VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn7 VSS D net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn6 net3 E net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn5 net4 net6 net3 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn4 net4 net1 VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn9 VSS net3 net0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn8 net0 SETN net1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3_56 net5 net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3 net5 net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn0 Q net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn0_11 Q net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn0_12 Q net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn0_11_1 Q net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp2 net6 E VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp6 VDD D net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net7 net6 net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 net3 E net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net8 net1 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 VDD net3 net1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp8 net1 SETN VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp7_53 net5 net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp7 net5 net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp0 Q net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp0_8 Q net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp0_32 Q net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp0_8_30 Q net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   MUX2_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:48:13 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT MUX2_X1 I0 I1 S Z VDD VNW VPW VSS 
*.PININFO I0:I I1:I S:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=((S * I1) + (!S * I0))
M_MN2 VSS int04 Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_MN4 net_1 I1 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_MN8 int04 S net_1 VPW nmos_5p0 W=0.660000U L=0.600000U
M_MN7 net_3 sel1_n int04 VPW nmos_5p0 W=0.660000U L=0.600000U
M_MN3 VSS I0 net_3 VPW nmos_5p0 W=0.660000U L=0.600000U
M_MN1 sel1_n S VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_MP5 VDD int04 Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_MP4 net_0 I1 VDD VNW pmos_5p0 W=0.915000U L=0.500000U
M_MP8 int04 sel1_n net_0 VNW pmos_5p0 W=0.915000U L=0.500000U
M_MP7 net_2 S int04 VNW pmos_5p0 W=0.915000U L=0.500000U
M_MP3 VDD I0 net_2 VNW pmos_5p0 W=0.915000U L=0.500000U
M_MP1 sel1_n S VDD VNW pmos_5p0 W=0.915000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   MUX2_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:48:10 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT MUX2_X2 I0 I1 S Z VDD VNW VPW VSS 
*.PININFO I0:I I1:I S:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=((S * I1) + (!S * I0))
M_MN2_12 VSS int04 Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_MN2 VSS int04 Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_MN4 net_1 I1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_MN8 int04 S net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_MN7 net_3 sel1_n int04 VPW nmos_5p0 W=1.320000U L=0.600000U
M_MN3 VSS I0 net_3 VPW nmos_5p0 W=1.320000U L=0.600000U
M_MN1 sel1_n S VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_MP5_6 VDD int04 Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_MP5 VDD int04 Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_MP4 net_0 I1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_MP8 int04 sel1_n net_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_MP7 net_2 S int04 VNW pmos_5p0 W=1.830000U L=0.500000U
M_MP3 VDD I0 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_MP1 sel1_n S VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   MUX2_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:48:11 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT MUX2_X4 I0 I1 S Z VDD VNW VPW VSS 
*.PININFO I0:I I1:I S:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=((S * I1) + (!S * I0))
M_MN2_12_7 VSS int04 Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_MN2_8 VSS int04 Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_MN2_12 VSS int04 Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_MN2 VSS int04 Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_MN4 net_1 I1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_MN8 int04 S net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_MN7 net_3 sel1_n int04 VPW nmos_5p0 W=1.320000U L=0.600000U
M_MN3 VSS I0 net_3 VPW nmos_5p0 W=1.320000U L=0.600000U
M_MN1 sel1_n S VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_MP5_6_5 VDD int04 Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_MP5_0 VDD int04 Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_MP5_6 VDD int04 Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_MP5 VDD int04 Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_MP4 net_0 I1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_MP8 int04 sel1_n net_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_MP7 net_2 S int04 VNW pmos_5p0 W=1.830000U L=0.500000U
M_MP3 VDD I0 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_MP1 sel1_n S VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   MUX4_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:47:43 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT MUX4_X1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS 
*.PININFO I0:I I1:I I2:I I3:I S0:I S1:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=((S0 * ((S1 * I3) + (!S1 * I1))) + (!S0 * ((S1 * I2) + (!S1 * I0))))
M_MN5 int01 I2 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_MN9 int02 sel1_n int01 VPW nmos_5p0 W=0.660000U L=0.600000U
M_MN10 int07 S0 int02 VPW nmos_5p0 W=0.660000U L=0.600000U
M_MN6 VSS I3 int07 VPW nmos_5p0 W=0.660000U L=0.600000U
M_instance_22 Z int03 VSS VPW nmos_5p0 W=0.900000U L=0.600000U
M_MN12 int03 S1 int02 VPW nmos_5p0 W=0.660000U L=0.600000U
M_MN11 int04 sel2_n int03 VPW nmos_5p0 W=0.660000U L=0.600000U
M_MN2 VSS S1 sel2_n VPW nmos_5p0 W=0.660000U L=0.600000U
M_MN4 int06 I1 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_MN8 int04 S0 int06 VPW nmos_5p0 W=0.660000U L=0.600000U
M_MN7 int05 sel1_n int04 VPW nmos_5p0 W=0.660000U L=0.600000U
M_MN3 VSS I0 int05 VPW nmos_5p0 W=0.660000U L=0.600000U
M_MN1 sel1_n S0 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_MP2 int01 I2 VDD VNW pmos_5p0 W=0.915000U L=0.500000U
M_MP9 int02 S0 int01 VNW pmos_5p0 W=0.915000U L=0.500000U
M_MP10 int07 sel1_n int02 VNW pmos_5p0 W=0.915000U L=0.500000U
M_MP6 VDD I3 int07 VNW pmos_5p0 W=0.915000U L=0.500000U
M_instance_1 Z int03 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_MP12 int03 sel2_n int02 VNW pmos_5p0 W=0.915000U L=0.500000U
M_MP11 int04 S1 int03 VNW pmos_5p0 W=0.915000U L=0.500000U
M_MP5 VDD S1 sel2_n VNW pmos_5p0 W=0.915000U L=0.500000U
M_MP4 int06 I1 VDD VNW pmos_5p0 W=0.915000U L=0.500000U
M_MP8 int04 sel1_n int06 VNW pmos_5p0 W=0.915000U L=0.500000U
M_MP7 int05 S0 int04 VNW pmos_5p0 W=0.915000U L=0.500000U
M_MP3 VDD I0 int05 VNW pmos_5p0 W=0.915000U L=0.500000U
M_MP1 sel1_n S0 VDD VNW pmos_5p0 W=0.915000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   MUX4_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs008             *
* at 11:47:41 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT MUX4_X2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS 
*.PININFO I0:I I1:I I2:I I3:I S0:I S1:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=((S0 * ((S1 * I3) + (!S1 * I1))) + (!S0 * ((S1 * I2) + (!S1 * I0))))
M_MN5 int01 I2 VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN9 int02 sel1_n int01 VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN10 int07 S0 int02 VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN6 VSS I3 int07 VPW nmos_5p0 W=0.800000U L=0.600000U
M_instance_22 Z int03 VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_instance_22_11 Z int03 VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN12 int03 S1 int02 VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN11 int04 sel2_n int03 VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN2 VSS S1 sel2_n VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN4 int06 I1 VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN8 int04 S0 int06 VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN7 int05 sel1_n int04 VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN3 VSS I0 int05 VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN1 sel1_n S0 VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_MP2 int01 I2 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP9 int02 S0 int01 VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP10 int07 sel1_n int02 VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP6 VDD I3 int07 VNW pmos_5p0 W=1.280000U L=0.500000U
M_instance_1 Z int03 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_instance_1_6 Z int03 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP12 int03 sel2_n int02 VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP11 int04 S1 int03 VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP5 VDD S1 sel2_n VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP4 int06 I1 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP8 int04 sel1_n int06 VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP7 int05 S0 int04 VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP3 VDD I0 int05 VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP1 sel1_n S0 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   MUX4_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs008             *
* at 11:47:40 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT MUX4_X4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS 
*.PININFO I0:I I1:I I2:I I3:I S0:I S1:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=((S0 * ((S1 * I3) + (!S1 * I1))) + (!S0 * ((S1 * I2) + (!S1 * I0))))
M_MN5 int01 I2 VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN9 int02 sel1_n int01 VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN10 int07 S0 int02 VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN6 VSS I3 int07 VPW nmos_5p0 W=0.800000U L=0.600000U
M_instance_22 Z int03 VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_instance_22_11 Z int03 VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_instance_22_18 Z int03 VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_instance_22_11_19 Z int03 VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN12 int03 S1 int02 VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN11 int04 sel2_n int03 VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN2 VSS S1 sel2_n VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN4 int06 I1 VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN8 int04 S0 int06 VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN7 int05 sel1_n int04 VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN3 VSS I0 int05 VPW nmos_5p0 W=0.800000U L=0.600000U
M_MN1 sel1_n S0 VSS VPW nmos_5p0 W=0.800000U L=0.600000U
M_MP2 int01 I2 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP9 int02 S0 int01 VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP10 int07 sel1_n int02 VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP6 VDD I3 int07 VNW pmos_5p0 W=1.280000U L=0.500000U
M_instance_1 Z int03 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_instance_1_6 Z int03 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_instance_1_9 Z int03 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_instance_1_6_3 Z int03 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP12 int03 sel2_n int02 VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP11 int04 S1 int03 VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP5 VDD S1 sel2_n VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP4 int06 I1 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP8 int04 sel1_n int06 VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP7 int05 S0 int04 VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP3 VDD I0 int05 VNW pmos_5p0 W=1.280000U L=0.500000U
M_MP1 sel1_n S0 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NAND2_X1.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:48:24 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT NAND2_X1 A1 A2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(A1 * A2)
M_i_1 net_0 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 ZN A2 VDD VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_2 VDD A1 ZN VNW pmos_5p0 W=1.645000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NAND2_X2.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:48:26 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT NAND2_X2 A1 A2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(A1 * A2)
M_i_1_1 net_0_0 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 ZN A1 net_0_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 net_0_1 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 VSS A2 net_0_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 ZN A2 VDD VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_2_1 VDD A1 ZN VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_2_0 ZN A1 VDD VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_3_0 VDD A2 ZN VNW pmos_5p0 W=1.645000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NAND2_X4.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:29 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT NAND2_X4 A1 A2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(A1 * A2)
M_i_1_3 net_0_0 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 ZN A1 net_0_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 net_0_1 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_2 VSS A2 net_0_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 net_0_2 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 ZN A1 net_0_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 net_0_3 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 VSS A2 net_0_3 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_3 ZN A2 VDD VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_2_3 VDD A1 ZN VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_2_2 ZN A1 VDD VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_3_2 VDD A2 ZN VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_3_1 ZN A2 VDD VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_2_1 VDD A1 ZN VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_2_0 ZN A1 VDD VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_3_0 VDD A2 ZN VNW pmos_5p0 W=1.645000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NAND3_X1.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs024             *
* at 11:48:09 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT NAND3_X1 A1 A2 A3 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!((A1 * A2) * A3)
M_i_2 net_1 A3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1 net_0 A2 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5 ZN A3 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_4 VDD A2 ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_3 ZN A1 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NAND3_X2.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:48:06 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT NAND3_X2 A1 A2 A3 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!((A1 * A2) * A3)
M_i_2_1 net_1_0 A3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 net_0_0 A2 net_1_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 ZN A1 net_0_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 net_0_1 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 net_1_1 A2 net_0_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 VSS A3 net_1_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_1 ZN A3 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_4_0 VDD A2 ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_3_0 ZN A1 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_3_1 VDD A1 ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_4_1 ZN A2 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_5_0 VDD A3 ZN VNW pmos_5p0 W=1.460000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NAND3_X4.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs010             *
* at 11:48:06 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT NAND3_X4 A1 A2 A3 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!((A1 * A2) * A3)
M_i_1_3 net_1_3 A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 VSS A3 net_1_3 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 net_1_2 A3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_2 net_0 A2 net_1_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 net_1_1 A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_2 VSS A3 net_1_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_3 net_1_0 A3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 net_0_0 A2 net_1_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 ZN A1 net_0_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_3 ZN A2 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_5_0 VDD A3 ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_5_1 ZN A3 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_4_2 VDD A2 ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_4_1 ZN A2 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_5_2 VDD A3 ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_5_3 ZN A3 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_4_0 VDD A2 ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_3_3 ZN A1 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_3_2 VDD A1 ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_3_1 ZN A1 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_3_0 VDD A1 ZN VNW pmos_5p0 W=1.460000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NAND4_X1.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs007             *
* at 11:47:59 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT NAND4_X1 A1 A2 A3 A4 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 * A2) * A3) * A4)
M_i_3 net_2 A4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2 net_1 A3 net_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1 net_0 A2 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_7 ZN A4 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_6 VDD A3 ZN VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_5 ZN A2 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_4 VDD A1 ZN VNW pmos_5p0 W=1.280000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NAND4_X2.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:47:59 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT NAND4_X2 A1 A2 A3 A4 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 * A2) * A3) * A4)
M_i_3_0 net_2_0 A4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_1_0 A3 net_2_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 net_0_0 A2 net_1_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 ZN A1 net_0_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 net_0_1 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 net_1_1 A2 net_0_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 net_2_1 A3 net_1_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 VSS A4 net_2_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_7_0 VDD A4 ZN VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_6_0 ZN A3 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_5_0 VDD A2 ZN VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_4_0 ZN A1 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_4_1 VDD A1 ZN VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_5_1 ZN A2 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_6_1 VDD A3 ZN VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_7_1 ZN A4 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NAND4_X4.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs021             *
* at 11:48:03 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT NAND4_X4 A1 A2 A3 A4 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 * A2) * A3) * A4)
M_i_2_3 net_2_3 A3 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_3 VSS A4 net_2_3 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_2 net_2_2 A4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_2 net_1 A3 net_2_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 net_2_1 A3 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 VSS A4 net_2_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 net_2_0 A4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_1_0 A3 net_2_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_3 net_0_3 A2 net_1_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 ZN A1 net_0_3 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 net_0_2 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_2 net_1 A2 net_0_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 net_0_1 A2 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 ZN A1 net_0_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 net_0_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 net_1 A2 net_0_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_3 ZN A3 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_7_3 VDD A4 ZN VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_7_2 ZN A4 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_6_2 VDD A3 ZN VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_6_1 ZN A3 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_7_1 VDD A4 ZN VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_7_0 ZN A4 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_6_0 VDD A3 ZN VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_5_3 ZN A2 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_4_3 VDD A1 ZN VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_4_2 ZN A1 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_5_2 VDD A2 ZN VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_5_1 ZN A2 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_4_1 VDD A1 ZN VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_4_0 ZN A1 VDD VNW pmos_5p0 W=1.280000U L=0.500000U
M_i_5_0 VDD A2 ZN VNW pmos_5p0 W=1.280000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NOR2_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:24 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT NOR2_X1 A1 A2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(A1 + A2)
M_i_1 ZN A2 VSS VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_0 VSS A1 ZN VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_3 net_0 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_2 ZN A1 net_0 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NOR2_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:26 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT NOR2_X2 A1 A2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(A1 + A2)
M_i_1_1 ZN A2 VSS VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_0_1 VSS A1 ZN VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_0_0 ZN A1 VSS VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_1_0 VSS A2 ZN VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_3_1 net_0_0 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_2_1 ZN A1 net_0_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_2_0 net_0_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0 VDD A2 net_0_1 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NOR2_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:27 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT NOR2_X4 A1 A2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(A1 + A2)
M_i_1_3 ZN A2 VSS VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_0_3 VSS A1 ZN VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_0_2 ZN A1 VSS VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_1_2 VSS A2 ZN VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_1_1 ZN A2 VSS VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_0_1 VSS A1 ZN VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_0_0 ZN A1 VSS VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_1_0 VSS A2 ZN VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_3_3 net_0_0 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_2_3 ZN A1 net_0_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_2_2 net_0_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_2 VDD A2 net_0_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 net_0_2 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_2_1 ZN A1 net_0_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_2_0 net_0_3 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0 VDD A2 net_0_3 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NOR3_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs027             *
* at 11:48:01 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT NOR3_X1 A1 A2 A3 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!((A1 + A2) + A3)
M_i_2 ZN A3 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_1 VSS A2 ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_0 ZN A1 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_5 net_1 A3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4 net_0 A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3 ZN A1 net_0 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NOR3_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:48:03 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT NOR3_X2 A1 A2 A3 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!((A1 + A2) + A3)
M_i_2_1 VSS A3 ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_1_0 ZN A2 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_0_0 VSS A1 ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_0_1 ZN A1 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_1_1 VSS A2 ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_2_0 ZN A3 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_5_1 net_1_0 A3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 net_0_0 A2 net_1_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0 ZN A1 net_0_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 net_0_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 net_1_1 A2 net_0_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 VDD A3 net_1_1 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NOR3_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:48:04 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT NOR3_X4 A1 A2 A3 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!((A1 + A2) + A3)
M_i_1_3 ZN A2 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_2_0 VSS A3 ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_2_1 ZN A3 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_1_2 VSS A2 ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_1_1 ZN A2 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_2_2 VSS A3 ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_2_3 ZN A3 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_1_0 VSS A2 ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_0_3 ZN A1 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_0_2 VSS A1 ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_0_1 ZN A1 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_0_0 VSS A1 ZN VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_4_3 net_1_3 A2 net_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 VDD A3 net_1_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 net_1_2 A3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_2 net_0 A2 net_1_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 net_1_1 A2 net_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_2 VDD A3 net_1_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_3 net_1_0 A3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 net_0_0 A2 net_1_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_3 ZN A1 net_0_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_2 net_0 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 ZN A1 net_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0 net_0 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NOR4_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:47:57 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT NOR4_X1 A1 A2 A3 A4 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) + A3) + A4)
M_i_3 ZN A4 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_2 VSS A3 ZN VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_1 ZN A2 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_0 VSS A1 ZN VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_7 net_2 A4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 net_1 A3 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5 net_0 A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4 ZN A1 net_0 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NOR4_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:47:59 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT NOR4_X2 A1 A2 A3 A4 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) + A3) + A4)
M_i_2_1 ZN A3 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_3_1 VSS A4 ZN VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_3_0 ZN A4 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_2_0 VSS A3 ZN VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_1_1 ZN A2 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_0_1 VSS A1 ZN VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_0_0 ZN A1 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_1_0 VSS A2 ZN VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_6_1 net_2_1 A3 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 VDD A4 net_2_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 net_2_0 A4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 net_1_0 A3 net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 net_0_1 A2 net_1_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 ZN A1 net_0_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 net_0_0 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 net_1 A2 net_0_0 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   NOR4_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:47:56 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT NOR4_X4 A1 A2 A3 A4 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) + A3) + A4)
M_i_2_3 ZN A3 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_3_3 VSS A4 ZN VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_3_2 ZN A4 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_2_2 VSS A3 ZN VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_2_1 ZN A3 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_3_1 VSS A4 ZN VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_3_0 ZN A4 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_2_0 VSS A3 ZN VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_1_3 ZN A2 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_0_3 VSS A1 ZN VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_0_2 ZN A1 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_1_2 VSS A2 ZN VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_1_1 ZN A2 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_0_1 VSS A1 ZN VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_0_0 ZN A1 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_1_0 VSS A2 ZN VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_6_3 net_2_3 A3 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_3 VDD A4 net_2_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_2 net_2_2 A4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_2 net_1 A3 net_2_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 net_2_1 A3 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 VDD A4 net_2_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 net_2_0 A4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 net_1_0 A3 net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_3 net_0_3 A2 net_1_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_3 ZN A1 net_0_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_2 net_0_2 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_2 net_1 A2 net_0_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 net_0_1 A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 ZN A1 net_0_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 net_0_0 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 net_1 A2 net_0_0 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI211_X1.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:47:47 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI211_X1 A1 A2 B C ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B:I C:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) * B) * C)
M_i_1 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2 net_1 B net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 VSS C net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5 net_2 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4 ZN A1 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 VDD B ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_7 ZN C VDD VNW pmos_5p0 W=1.460000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI211_X2.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:47:48 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI211_X2 A1 A2 B C ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B:I C:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) * B) * C)
M_i_1_1 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_1_0 B net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 VSS C net_1_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 net_1_1 C VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 net_0 B net_1_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_1 net_2_0 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 ZN A1 net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 net_2_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 VDD A2 net_2_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 ZN B VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_7_0 VDD C ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_7_1 ZN C VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_6_1 VDD B ZN VNW pmos_5p0 W=1.460000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI211_X4.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs016             *
* at 11:47:50 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI211_X4 A1 A2 B C ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B:I C:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) * B) * C)
M_i_1_3 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_2 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_1_0 B net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 VSS C net_1_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 net_1_1 C VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 net_0 B net_1_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_2 net_1_2 B net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_2 VSS C net_1_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_3 net_1_3 C VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_3 net_0 B net_1_3 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_3 net_2_0 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_3 ZN A1 net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_2 net_2_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_2 VDD A2 net_2_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 net_2_2 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 ZN A1 net_2_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 net_2_3 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 VDD A2 net_2_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 ZN B VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_7_0 VDD C ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_7_1 ZN C VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_6_1 VDD B ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_6_2 ZN B VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_7_2 VDD C ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_7_3 ZN C VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_6_3 VDD B ZN VNW pmos_5p0 W=1.460000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI21_X1.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:03 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI21_X1 A1 A2 B ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!((A1 + A2) * B)
M_i_1 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2 VSS B net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4 net_1 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3 ZN A1 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5 VDD B ZN VNW pmos_5p0 W=1.645000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI21_X2.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:03 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI21_X2 A1 A2 B ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!((A1 + A2) * B)
M_i_2_1 VSS B net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_0 B VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_1 ZN B VDD VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_5_0 VDD B ZN VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_4_1 net_1_0 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 ZN A1 net_1_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0 net_1_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 VDD A2 net_1_1 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI21_X4.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:07 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI21_X4 A1 A2 B ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!((A1 + A2) * B)
M_i_1_3 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_2 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_3 VSS B net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_2 net_0 B VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 VSS B net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_0 B VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_3 net_1_0 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_3 ZN A1 net_1_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_2 net_1_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_2 VDD A2 net_1_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 net_1_2 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 ZN A1 net_1_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0 net_1_3 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 VDD A2 net_1_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_3 ZN B VDD VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_5_2 VDD B ZN VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_5_1 ZN B VDD VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_5_0 VDD B ZN VNW pmos_5p0 W=1.645000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI221_X1.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:47:41 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI221_X1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B1:I B2:I C:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) * (B1 + B2)) * C)
M_i_4 VSS B2 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 net_1 B1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2 net_0 C net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_9 net_3 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8 ZN B1 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7 VDD C ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_6 net_2 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5 ZN A1 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI221_X2.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs027             *
* at 11:47:41 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI221_X2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B1:I B2:I C:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) * (B1 + B2)) * C)
M_i_2_1 net_1 C net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_1 VSS B2 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 net_1 B1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 VSS B1 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_0 net_1 B2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_0 C net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_7_1 VDD C ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_9_1 net_3_0 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_1 ZN B1 net_3_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_0 net_3_1 B1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_0 VDD B2 net_3_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 ZN C VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_5_1 net_2_0 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 VDD A2 net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 net_2_1 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 ZN A1 net_2_1 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI221_X4.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:47:47 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI221_X4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B1:I B2:I C:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) * (B1 + B2)) * C)
M_i_3_3 net_1 B1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_3 VSS B2 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_2 net_1 B2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_2 VSS B1 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 net_1 B1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_1 VSS B2 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_0 net_1 B2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 VSS B1 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_3 net_1 C net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_2 net_0 C net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 net_1 C net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_0 C net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_3 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_2 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_8_3 net_3_0 B1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_3 VDD B2 net_3_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_2 net_3_1 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_2 ZN B1 net_3_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_1 net_3_2 B1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_1 VDD B2 net_3_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_0 net_3_3 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_0 ZN B1 net_3_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_3 VDD C ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_7_2 ZN C VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_7_1 VDD C ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_7_0 ZN C VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_5_3 net_2_0 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_3 VDD A2 net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_2 net_2_1 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_2 ZN A1 net_2_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 net_2_2 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 VDD A2 net_2_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 net_2_3 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 ZN A1 net_2_3 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI222_X1.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:47:24 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI222_X1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) * (B1 + B2)) * (C1 + C2))
M_i_5 net_1 C2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4 VSS C1 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2 net_1 B1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 net_0 B2 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_11 net_4 C2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10 ZN C1 net_4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8 net_3 B1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9 VDD B2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7 net_2 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 ZN A1 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI222_X2.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:47:22 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI222_X2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) * (B1 + B2)) * (C1 + C2))
M_i_4_1 net_1 C1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_1 VSS C2 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_0 net_1 C2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_0 VSS C1 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_1 B1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 net_0 B2 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 net_1 B2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 net_0 B1 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_10_1 net_4_1 C1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_1 VDD C2 net_4_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_0 net_4_0 C2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10_0 ZN C1 net_4_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_0 net_3_1 B1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_0 VDD B2 net_3_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_1 net_3_0 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_1 ZN B1 net_3_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 net_2_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 VDD A2 net_2_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 net_2_0 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 ZN A1 net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI222_X4.                                                       *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:47:28 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI222_X4 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) * (B1 + B2)) * (C1 + C2))
M_i_4_3 net_1 C1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_3 VSS C2 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_2 net_1 C2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_2 VSS C1 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_1 net_1 C1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_1 VSS C2 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_0 net_1 C2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_0 VSS C1 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_1 B1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 net_0 B2 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 net_1 B2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 net_0 B1 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_2 net_1 B1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_2 net_0 B2 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_3 net_1 B2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_3 net_0 B1 net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_2 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_3 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_10_3 net_4_3 C1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_3 VDD C2 net_4_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_2 net_4_2 C2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10_2 ZN C1 net_4_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10_1 net_4_1 C1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_1 VDD C2 net_4_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_0 net_4_0 C2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10_0 ZN C1 net_4_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_0 net_3_3 B1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_0 VDD B2 net_3_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_1 net_3_2 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_1 ZN B1 net_3_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_2 net_3_1 B1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_2 VDD B2 net_3_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_3 net_3_0 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_3 ZN B1 net_3_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 net_2_3 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 VDD A2 net_2_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 net_2_2 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 ZN A1 net_2_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_2 net_2_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_2 VDD A2 net_2_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_3 net_2_0 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_3 ZN A1 net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI22_X1.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:47:52 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI22_X1 A1 A2 B1 B2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B1:I B2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!((A1 + A2) * (B1 + B2))
M_i_3 VSS B2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2 net_0 B1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_7 net_2 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 ZN B1 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4 net_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5 VDD A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI22_X2.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs024             *
* at 11:47:54 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI22_X2 A1 A2 B1 B2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B1:I B2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!((A1 + A2) * (B1 + B2))
M_i_3_1 VSS B2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 net_0 B1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 VSS B1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 net_0 B2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_7_1 net_2_0 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 ZN B1 net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 net_2_1 B1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 VDD B2 net_2_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 net_1_0 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 ZN A1 net_1_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 net_1_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 VDD A2 net_1_1 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI22_X4.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:47:56 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI22_X4 A1 A2 B1 B2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I B1:I B2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!((A1 + A2) * (B1 + B2))
M_i_3_3 VSS B2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_3 net_0 B1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_2 VSS B1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_2 net_0 B2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 VSS B2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 net_0 B1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 VSS B1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 net_0 B2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_2 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_3 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_7_3 net_2_0 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_3 ZN B1 net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_2 net_2_1 B1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_2 VDD B2 net_2_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 net_2_2 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 ZN B1 net_2_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 net_2_3 B1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 VDD B2 net_2_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 net_1_0 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 ZN A1 net_1_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 net_1_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 VDD A2 net_1_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_2 net_1_2 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_2 ZN A1 net_1_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_3 net_1_3 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_3 VDD A2 net_1_3 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI31_X1.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs024             *
* at 11:47:50 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI31_X1 A1 A2 A3 B ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I B:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) + A3) * B)
M_i_3 net_0 B VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2 ZN A3 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_7 ZN B VDD VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_4 net_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5 net_2 A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 VDD A3 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI31_X2.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:47:48 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI31_X2 A1 A2 A3 B ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I B:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) + A3) * B)
M_i_3_1 VSS B net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 net_0 B VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 ZN A3 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_0 A3 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_7_1 ZN B VDD VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_7_0 VDD B ZN VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_6_1 net_2_0 A3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 net_1_0 A2 net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 ZN A1 net_1_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 net_1_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 net_2_1 A2 net_1_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 VDD A3 net_2_1 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI31_X4.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:47:53 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI31_X4 A1 A2 A3 B ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I B:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) + A3) * B)
M_i_2_3 ZN A3 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_2 net_0 A3 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 ZN A3 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_0 A3 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_3 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_2 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_3 VSS B net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_2 net_0 B VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 VSS B net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 net_0 B VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_3 VDD A3 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_2 net_2 A3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 VDD A3 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 net_2_0 A3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_3 net_1_0 A2 net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_3 ZN A1 net_1_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_2 net_1_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_2 net_2 A2 net_1_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 net_1_2 A2 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 ZN A1 net_1_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 net_1_3 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 net_2 A2 net_1_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_3 ZN B VDD VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_7_2 VDD B ZN VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_7_1 ZN B VDD VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_7_0 VDD B ZN VNW pmos_5p0 W=1.645000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI32_X1.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs021             *
* at 11:47:42 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI32_X1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I B1:I B2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) + A3) * (B1 + B2))
M_i_4 net_0 A3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 VSS A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2 net_0 A1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0 ZN B1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1 net_0 B2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_9 net_3 A3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8 net_2 A2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7 ZN A1 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5 net_1 B1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 VDD B2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI32_X2.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:47:42 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI32_X2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I B1:I B2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) + A3) * (B1 + B2))
M_i_4_1 VSS A3 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 net_0 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 VSS A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_0 A1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 VSS A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_0 net_0 A3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 ZN B2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 net_0 B1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 ZN B1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 net_0 B2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_9_1 net_3_0 A3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_1 net_2_0 A2 net_3_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 ZN A1 net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 net_2_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_0 net_3_1 A2 net_2_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_0 VDD A3 net_3_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 net_1_0 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 ZN B1 net_1_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 net_1_1 B1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 VDD B2 net_1_1 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI32_X4.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:47:46 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI32_X4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I B1:I B2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) + A3) * (B1 + B2))
M_i_3_3 VSS A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_3 net_0 A3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_2 VSS A3 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_2 net_0 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 VSS A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_1 net_0 A3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_0 VSS A3 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 net_0 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_3 VSS A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_2 net_0 A1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 VSS A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 net_0 A1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_3 ZN B2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 net_0 B1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 ZN B1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_2 net_0 B2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 ZN B2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 net_0 B1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 ZN B1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 net_0 B2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_8_3 net_3_0 A2 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_3 VDD A3 net_3_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_2 net_3_1 A3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_2 net_2 A2 net_3_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_1 net_3_2 A2 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_1 VDD A3 net_3_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_0 net_3_3 A3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_0 net_2_0 A2 net_3_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_3 ZN A1 net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_2 net_2 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 ZN A1 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 net_2 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_3 net_1_0 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_3 ZN B1 net_1_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_2 net_1_1 B1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_2 VDD B2 net_1_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 net_1_2 B2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 ZN B1 net_1_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 net_1_3 B1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 VDD B2 net_1_3 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI33_X1.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:47:28 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI33_X1 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) + A3) * ((B1 + B2) + B3))
M_i_5 net_0 B3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4 VSS B2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 net_0 B1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2 ZN A3 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_11 net_4 B3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10 net_3 B2 net_4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9 ZN B1 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 net_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7 net_2 A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8 VDD A3 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI33_X2.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:47:29 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI33_X2 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) + A3) * ((B1 + B2) + B3))
M_i_5_0 VSS B3 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_1 net_0 B2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 VSS B1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 net_0 B1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_0 VSS B2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_1 net_0 B3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 ZN A3 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 net_0 A3 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_11_0 net_4_0 B3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10_1 net_3_0 B2 net_4_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_1 ZN B1 net_3_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_0 net_3_1 B1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10_0 net_4_1 B2 net_3_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_1 VDD B3 net_4_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_0 net_2_0 A3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 net_1_0 A2 net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 ZN A1 net_1_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 net_1_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 net_2_1 A2 net_1_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_1 VDD A3 net_2_1 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OAI33_X4.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:47:37 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OAI33_X4 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(((A1 + A2) + A3) * ((B1 + B2) + B3))
M_i_4_0 VSS B2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_0 net_0 B3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_1 VSS B3 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_1 net_0 B2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_2 VSS B2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_2 net_0 B3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_3 VSS B3 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_3 net_0 B2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 VSS B1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 net_0 B1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_2 VSS B1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_3 net_0 B1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_3 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_3 net_0 A3 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_2 ZN A3 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_2 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 net_0 A3 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 ZN A3 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_10_0 net_4_0 B2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_0 VDD B3 net_4_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_1 net_4_1 B3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10_1 net_3 B2 net_4_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10_2 net_4_2 B2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_2 VDD B3 net_4_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_3 net_4_3 B3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10_3 net_3_0 B2 net_4_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_0 ZN B1 net_3_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_1 net_3 B1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_2 ZN B1 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_3 net_3 B1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 ZN A1 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 net_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_2 ZN A1 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_3 net_1_0 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_3 net_2_0 A2 net_1_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_3 VDD A3 net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_2 net_2_1 A3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_2 net_1 A2 net_2_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 net_2_2 A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_1 VDD A3 net_2_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_0 net_2_3 A3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 net_1 A2 net_2_3 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OR2_X1.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:48:20 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OR2_X1 A1 A2 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=(A1 + A2)
M_i_2 Z_neg A1 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_3 VSS A2 Z_neg VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4 net_0 A1 Z_neg VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_5 VDD A2 net_0 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_1 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OR2_X2.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:48:21 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OR2_X2 A1 A2 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=(A1 + A2)
M_i_2 Z_neg A1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 VSS A2 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4 net_0 A1 Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5 VDD A2 net_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OR2_X4.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:48:24 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OR2_X4 A1 A2 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=(A1 + A2)
M_i_3_1 Z_neg A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 VSS A1 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 Z_neg A1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 VSS A2 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_1 net_0_1 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 Z_neg A1 net_0_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 net_0_0 A1 Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 VDD A2 net_0_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OR3_X1.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:04 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OR3_X1 A1 A2 A3 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=((A1 + A2) + A3)
M_i_2 VSS A1 Z_neg VPW nmos_5p0 W=0.525000U L=0.600000U
M_i_3 Z_neg A2 VSS VPW nmos_5p0 W=0.525000U L=0.600000U
M_i_4 VSS A3 Z_neg VPW nmos_5p0 W=0.525000U L=0.600000U
M_i_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5 net_0 A1 Z_neg VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_6 net_1 A2 net_0 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_7 VDD A3 net_1 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_1 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OR3_X2.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:02 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OR3_X2 A1 A2 A3 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=((A1 + A2) + A3)
M_i_2 VSS A1 Z_neg VPW nmos_5p0 W=1.050000U L=0.600000U
M_i_3 Z_neg A2 VSS VPW nmos_5p0 W=1.050000U L=0.600000U
M_i_4 VSS A3 Z_neg VPW nmos_5p0 W=1.050000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5 net_0 A1 Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 net_1 A2 net_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7 VDD A3 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OR3_X4.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:04 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OR3_X4 A1 A2 A3 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=((A1 + A2) + A3)
M_i_4_0 Z_neg A3 VSS VPW nmos_5p0 W=1.050000U L=0.600000U
M_i_3_1 VSS A2 Z_neg VPW nmos_5p0 W=1.050000U L=0.600000U
M_i_2_1 Z_neg A1 VSS VPW nmos_5p0 W=1.050000U L=0.600000U
M_i_2_0 VSS A1 Z_neg VPW nmos_5p0 W=1.050000U L=0.600000U
M_i_3_0 Z_neg A2 VSS VPW nmos_5p0 W=1.050000U L=0.600000U
M_i_4_1 VSS A3 Z_neg VPW nmos_5p0 W=1.050000U L=0.600000U
M_i_0_3 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_7_0 net_1_1 A3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 net_0_1 A2 net_1_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 Z_neg A1 net_0_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 net_0_0 A1 Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 net_1_0 A2 net_0_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 VDD A3 net_1_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OR4_X1.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:47:44 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OR4_X1 A1 A2 A3 A4 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I A4:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=(((A1 + A2) + A3) + A4)
M_i_2 Z_neg A1 VSS VPW nmos_5p0 W=0.395000U L=0.600000U
M_i_3 VSS A2 Z_neg VPW nmos_5p0 W=0.395000U L=0.600000U
M_i_4 Z_neg A3 VSS VPW nmos_5p0 W=0.395000U L=0.600000U
M_i_5 VSS A4 Z_neg VPW nmos_5p0 W=0.395000U L=0.600000U
M_i_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6 net_0 A1 Z_neg VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_7 net_1 A2 net_0 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_8 net_2 A3 net_1 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_9 VDD A4 net_2 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_1 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OR4_X2.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs007             *
* at 11:47:42 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OR4_X2 A1 A2 A3 A4 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I A4:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=(((A1 + A2) + A3) + A4)
M_i_2 Z_neg A1 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_3 VSS A2 Z_neg VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_4 Z_neg A3 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_5 VSS A4 Z_neg VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6 net_0 A1 Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7 net_1 A2 net_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8 net_2 A3 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9 VDD A4 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   OR4_X4.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs007             *
* at 11:47:45 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT OR4_X4 A1 A2 A3 A4 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I A4:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=(((A1 + A2) + A3) + A4)
M_i_5_1_x2_1 Z_neg A4 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_4_1_x2_1 VSS A3 Z_neg VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_3_1_x2_1 Z_neg A2 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_2_1_x2_1 VSS A1 Z_neg VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_2_1_x2_0 Z_neg A1 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_3_1_x2_0 VSS A2 Z_neg VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_4_1_x2_0 Z_neg A3 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_5_1_x2_0 VSS A4 Z_neg VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_0_3_x4_3 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3_x4_2 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3_x4_1 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3_x4_0 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_9_0_m2_1 net_2_0_1 A4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_0_m2_1 net_1_0_1 A3 net_2_0_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0_m2_1 net_0_0_1 A2 net_1_0_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0_m2_1 Z_neg A1 net_0_0_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0_m2_0 net_0_0_0 A1 Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0_m2_0 net_1_0_0 A2 net_0_0_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_0_m2_0 net_2_0_0 A3 net_1_0_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_0_m2_0 VDD A4 net_2_0_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3_x4_3 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3_x4_2 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3_x4_1 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3_x4_0 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFFQ_X1.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:46:42 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT SDFFQ_X1 D SE SI CLK Q VDD VNW VPW VSS 
*.PININFO D:I SE:I SI:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn14 net8 SE VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn12 net12 SI VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn13 net12 SE net6 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn8 net6 net8 net9n VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn10 VSS D net9n VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn16 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn9 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn11 net6 ncki net5 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn0 net5 cki net11 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn1 VSS net10 net11 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn15 net10 net5 VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn2 net0 cki net10 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn3 net7 ncki net0 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn4 VSS net1 net7 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn5 net1 net0 VSS VPW nmos_5p0 W=0.750000U L=0.600000U
M_tn6 Q net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp14 net8 SE VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 net3 SI VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net2 net8 net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp8 net9p SE net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 VDD D net9p VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp9 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp11 net5 cki net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp0 net4 ncki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp1 VDD net10 net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp15 net10 net5 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net0 ncki net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net7_p cki net0 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 VDD net1 net7_p VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net1 net0 VDD VNW pmos_5p0 W=1.100000U L=0.500000U
M_tp4 Q net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFFQ_X2.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:46:42 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT SDFFQ_X2 D SE SI CLK Q VDD VNW VPW VSS 
*.PININFO D:I SE:I SI:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn14 net8 SE VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn12 net12 SI VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn13 net12 SE net6 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn8 net6 net8 net9n VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn10 VSS D net9n VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn16 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn9 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn11 net6 ncki net5 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn0 net5 cki net11 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn1 VSS net10 net11 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn15 net10 net5 VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn2 net0 cki net10 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn3 net7 ncki net0 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn4 VSS net1 net7 VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn5 net1 net0 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn6_6 Q net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn6 Q net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp14 net8 SE VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 net3 SI VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net2 net8 net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp8 net9p SE net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 VDD D net9p VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp9 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp11 net5 cki net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp0 net4 ncki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp1 VDD net10 net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp15 net10 net5 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net0 ncki net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net7_p cki net0 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 VDD net1 net7_p VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp3 net1 net0 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4_12 Q net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4 Q net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFFQ_X4.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:46:43 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT SDFFQ_X4 D SE SI CLK Q VDD VNW VPW VSS 
*.PININFO D:I SE:I SI:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn14 net8 SE VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn12 net12 SI VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn13 net12 SE net6 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn8 net6 net8 net9n VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn10 VSS D net9n VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn16 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn9 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn11 net6 ncki net5 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn0 net5 cki net11 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn1 VSS net10 net11 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn15 net10 net5 VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn2 net0 cki net10 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn3 net7 ncki net0 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn4 VSS net1 net7 VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn5 net1 net0 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn6_6_25 Q net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn6_5 Q net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn6_6 Q net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn6 Q net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp14 net8 SE VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 net3 SI VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net2 net8 net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp8 net9p SE net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 VDD D net9p VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp9 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp11 net5 cki net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp0 net4 ncki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp1 VDD net10 net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp15 net10 net5 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net0 ncki net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net7_p cki net0 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 VDD net1 net7_p VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp3 net1 net0 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4_12_24 Q net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4_16 Q net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4_12 Q net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4 Q net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFFRNQ_X1.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:46:43 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT SDFFRNQ_X1 D RN SE SI CLK Q VDD VNW VPW VSS 
*.PININFO D:I RN:I SE:I SI:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn17 net3 SE VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn7 VSS SI net13 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn6 net13 SE net10 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn11 net10 D net5 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn16 net5 net3 VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn10 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn13 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn15 net10 ncki net1 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn14 net1 cki net15 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn8 net12 net2 net15 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn9 VSS RN net12 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn18 VSS net1 net2 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn0 net8 cki net2 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn1 net11 ncki net8 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn12 net11 net4 VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn5 net0 RN VSS VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn4 net4 net8 net0 VPW nmos_5p0 W=0.580000U L=0.600000U
M_tn3 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp17 net3 SE VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 net7 SI VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 net6 net3 net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 net14 D net6 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp14 VDD SE net14 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp8 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp11 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp15 net1 cki net6 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net9 ncki net1 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 VDD net2 net9 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net9 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 VDD net1 net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 net2 ncki net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net8 cki net11 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net11 net4 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net4 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 VDD net8 net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp1 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFFRNQ_X2.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:46:43 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT SDFFRNQ_X2 D RN SE SI CLK Q VDD VNW VPW VSS 
*.PININFO D:I RN:I SE:I SI:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn17 net3 SE VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn7 VSS SI net13 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net13 SE net10 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn11 net10 D net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn16 net5 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn10 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn13 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn15 net10 ncki net1 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net1 cki net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn8 net12 net2 net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn9 VSS RN net12 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn18 VSS net1 net2 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn0 net8 cki net2 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 net11 ncki net8 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn12 net11 net4 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 net0 RN VSS VPW nmos_5p0 W=1.000000U L=0.600000U
M_tn4 net4 net8 net0 VPW nmos_5p0 W=1.000000U L=0.600000U
M_tn3_17 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp17 net3 SE VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 net7 SI VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 net6 net3 net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 net14 D net6 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp14 VDD SE net14 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp8 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp11 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp15 net1 cki net6 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net9 ncki net1 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 VDD net2 net9 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net9 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 VDD net1 net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 net2 ncki net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net8 cki net11 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net11 net4 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net4 RN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp4 VDD net8 net4 VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp1_16 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFFRNQ_X4.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs010             *
* at 11:46:36 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT SDFFRNQ_X4 D RN SE SI CLK Q VDD VNW VPW VSS 
*.PININFO D:I RN:I SE:I SI:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn17 net3 SE VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn7 VSS SI net13 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net13 SE net10 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn11 net10 D net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn16 net5 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn10 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn13 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn15 net10 ncki net1 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net1 cki net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn8 net12 net2 net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn9 VSS RN net12 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn18 VSS net1 net2 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn0 net8 cki net2 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 net11 ncki net8 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn12 net11 net4 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 net0 RN VSS VPW nmos_5p0 W=1.000000U L=0.600000U
M_tn4 net4 net8 net0 VPW nmos_5p0 W=1.000000U L=0.600000U
M_tn3_17_4 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3_27 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3_17 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp17 net3 SE VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 net7 SI VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 net6 net3 net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 net14 D net6 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp14 VDD SE net14 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp8 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp11 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp15 net1 cki net6 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net9 ncki net1 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 VDD net2 net9 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net9 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 VDD net1 net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 net2 ncki net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net8 cki net11 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net11 net4 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net4 RN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp4 VDD net8 net4 VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp1_16_17 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1_25 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1_16 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFFRSNQ_X1.                                                     *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs016             *
* at 11:46:35 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT SDFFRSNQ_X1 D RN SE SETN SI CLK Q VDD VNW VPW VSS 
*.PININFO D:I RN:I SE:I SETN:I SI:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn12 net9 SE VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn9 VSS SI net17 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn10 net17 SE net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn0 net14 D net8 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn11 net8 net9 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn2 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn8 net14 ncki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 net3 cki net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net15 net4 net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn7 VSS RN net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn3 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net5 cki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net7 ncki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 net1 SETN net7 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn16 VSS net6 net1 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn18 net2 RN VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn17 net6 net5 net2 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn19 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp12 net9 SE VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp11 net12 SI VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp8 net10 net9 net12 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp0 net11 D net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 VDD SE net11 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp1 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp2 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp10 net3 cki net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net13 ncki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net13 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 VDD net3 net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp20 net4 ncki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp19 net5 cki net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 net7 SETN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp14 net7 net6 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 net6 RN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp15 VDD net5 net6 VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp17 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFFRSNQ_X2.                                                     *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs007             *
* at 11:46:36 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT SDFFRSNQ_X2 D RN SE SETN SI CLK Q VDD VNW VPW VSS 
*.PININFO D:I RN:I SE:I SETN:I SI:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn12 net9 SE VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn9 VSS SI net17 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn10 net17 SE net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn0 net14 D net8 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn11 net8 net9 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn2 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn8 net14 ncki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 net3 cki net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net15 net4 net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn7 VSS RN net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn3 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net5 cki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net7 ncki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 net1 SETN net7 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn16 VSS net6 net1 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn18 net2 RN VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn17 net6 net5 net2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn19 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn19_14 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp12 net9 SE VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp11 net12 SI VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp8 net10 net9 net12 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp0 net11 D net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 VDD SE net11 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp1 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp2 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp10 net3 cki net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net13 ncki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net13 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 VDD net3 net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp20 net4 ncki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp19 net5 cki net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 net7 SETN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp14 net7 net6 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 net6 RN VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp15 VDD net5 net6 VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp17 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp17_7 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFFRSNQ_X4.                                                     *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs007             *
* at 11:46:37 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT SDFFRSNQ_X4 D RN SE SETN SI CLK Q VDD VNW VPW VSS 
*.PININFO D:I RN:I SE:I SETN:I SI:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn12 net9 SE VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn9 VSS SI net17 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn10 net17 SE net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn0 net14 D net8 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn11 net8 net9 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn2 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn8 net14 ncki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 net3 cki net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net15 net4 net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn7 VSS RN net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn3 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net5 cki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net7 ncki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 net1 SETN net7 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn16 VSS net6 net1 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn18 net2 RN VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn17 net6 net5 net2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn19 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn19_14 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn19_12 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn19_14_0 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp12 net9 SE VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp11 net12 SI VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp8 net10 net9 net12 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp0 net11 D net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 VDD SE net11 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp1 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp2 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp10 net3 cki net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net13 ncki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net13 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 VDD net3 net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp20 net4 ncki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp19 net5 cki net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 net7 SETN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp14 net7 net6 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 net6 RN VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp15 VDD net5 net6 VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp17 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp17_7 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp17_8 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp17_7_4 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFFSNQ_X1.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs008             *
* at 11:46:30 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT SDFFSNQ_X1 D SE SETN SI CLK Q VDD VNW VPW VSS 
*.PININFO D:I SE:I SETN:I SI:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn11 net9 SE VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn7 VSS SI net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn9 net15 SE net13 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn10 net13 D net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn8 net16 net9 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn3 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn0 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn6 net13 ncki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net3 cki net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 VSS net4 net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn2 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net5 cki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn12 net7 ncki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net1 SETN net7 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 VSS net6 net1 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn18 net6 net5 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn16 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp11 net9 SE VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net11 SI VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp1 net8 net9 net11 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp8 net12 D net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 VDD SE net12 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp0 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp9 net3 cki net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net10 ncki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net4 net3 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 net5 ncki net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp17 net7 cki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net7 SETN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 VDD net6 net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 net6 net5 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp14 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFFSNQ_X2.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs008             *
* at 11:46:31 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT SDFFSNQ_X2 D SE SETN SI CLK Q VDD VNW VPW VSS 
*.PININFO D:I SE:I SETN:I SI:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn11 net9 SE VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn7 VSS SI net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn9 net15 SE net13 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn10 net13 D net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn8 net16 net9 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn3 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn0 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn6 net13 ncki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net3 cki net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 VSS net4 net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn2 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net5 cki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn12 net7 ncki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net1 SETN net7 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 VSS net6 net1 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn18 net6 net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn16 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn16_8 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp11 net9 SE VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net11 SI VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp1 net8 net9 net11 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp8 net12 D net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 VDD SE net12 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp0 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp9 net3 cki net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net10 ncki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net4 net3 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 net5 ncki net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp17 net7 cki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net7 SETN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 VDD net6 net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 net6 net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp14 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp14_2 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   SDFFSNQ_X4.                                                      *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs027             *
* at 11:46:32 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT SDFFSNQ_X4 D SE SETN SI CLK Q VDD VNW VPW VSS 
*.PININFO D:I SE:I SETN:I SI:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G 
M_tn11 net9 SE VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn7 VSS SI net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn9 net15 SE net13 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn10 net13 D net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn8 net16 net9 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn3 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn0 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn6 net13 ncki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net3 cki net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 VSS net4 net14 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn2 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net5 cki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn12 net7 ncki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net1 SETN net7 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 VSS net6 net1 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn18 net6 net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn18_45 net6 net5 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn16 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn16_8 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn16_23 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn16_8_32 VSS net6 Q VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp11 net9 SE VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net11 SI VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp1 net8 net9 net11 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp8 net12 D net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 VDD SE net12 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp0 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp9 net3 cki net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net10 ncki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net4 net3 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 net5 ncki net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp17 net7 cki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net7 SETN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 VDD net6 net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 net6 net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp16_52 net6 net5 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp14 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp14_2 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp14_18 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp14_2_28 VDD net6 Q VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   TIEH.                                                            *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs001             *
* at 11:49:03 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT TIEH Z VDD VNW VPW VSS 
*.PININFO Z:O VDD:P VNW:P VPW:P VSS:G 
M_n_tran_1 VSS A A VPW nmos_5p0 W=0.660000U L=0.600000U
M_p_tran_2 VDD A Z VNW pmos_5p0 W=0.900000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   TIEL.                                                            *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs022             *
* at 11:49:05 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT TIEL ZN VDD VNW VPW VSS 
*.PININFO ZN:O VDD:P VNW:P VPW:P VSS:G 
M_n_tran_1 VSS A ZN VPW nmos_5p0 W=0.660000U L=0.600000U
M_transistor_0 VDD A A VNW pmos_5p0 W=0.900000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   XNOR2_X1.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:24 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT XNOR2_X1 A1 A2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(!((A1 * A2) + !(A1 + A2)))
M_i_6 net_2 A2 I VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_7 VSS A1 net_2 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_2 net_0 I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_8 I A2 VDD VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_9 VDD A1 I VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_5 ZN I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3 net_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4 VDD A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   XNOR2_X2.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs016             *
* at 11:48:22 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT XNOR2_X2 A1 A2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(!((A1 * A2) + !(A1 + A2)))
M_i_8 I A2 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_9 VSS A1 I VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_4 Z_neg I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2 net_0 A1 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 VSS A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 ZN Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS Z_neg ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_10 net_2 A2 I VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_11 VDD A1 net_2 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_7 net_1 I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5 Z_neg A1 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 net_1 A2 Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 ZN Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   XNOR2_X4.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs025             *
* at 11:48:22 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT XNOR2_X4 A1 A2 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(!((A1 * A2) + !(A1 + A2)))
M_i_8 I A2 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_9 VSS A1 I VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_4 Z_neg I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2 net_0 A1 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 VSS A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 ZN Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS Z_neg ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 ZN Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 VSS Z_neg ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_10 net_2 A2 I VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_11 VDD A1 net_2 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_7 net_1 I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5 Z_neg A1 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 net_1 A2 Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 ZN Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 ZN Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD Z_neg ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   XNOR3_X1.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:09 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT XNOR3_X1 A1 A2 A3 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(!((!((A1 * A2) + !(A1 + A2)) * A3) + !(!((A1 * A2) + !(A1 + A2)) + A3)))
M_i_12 I A2 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_13 VSS A1 I VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 I2 I VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_0 net_0 A1 I2 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_1 VSS A2 net_0 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_16 net_5 I2 I3 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_17 VSS A3 net_5 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_8 net_2 I3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6 ZN A3 net_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_7 net_2 I2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_14 net_4 A2 I VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_15 VDD A1 net_4 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_5 net_1 I VDD VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_3 I2 A1 net_1 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_4 net_1 A2 I2 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_18 I3 I2 VDD VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_19 VDD A3 I3 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_11 ZN I3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9 net_3 A3 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10 VDD I2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   XNOR3_X2.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:07 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT XNOR3_X2 A1 A2 A3 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(!((!((A1 * A2) + !(A1 + A2)) * A3) + !(!((A1 * A2) + !(A1 + A2)) + A3)))
M_i_14 I A2 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_15 VSS A1 I VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 I2 I VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_0 net_0 A1 I2 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_1 VSS A2 net_0 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_18 I3 I2 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_19 VSS A3 I3 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_10 Z_neg I3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_8 net_2 A3 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_9 VSS I2 net_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_1 VSS Z_neg ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_0 ZN Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_16 net_4 A2 I VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_17 VDD A1 net_4 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_5 net_1 I VDD VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_3 I2 A1 net_1 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_4 net_1 A2 I2 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_20 net_5 I2 I3 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_21 VDD A3 net_5 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_13 net_3 I3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11 Z_neg A3 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_12 net_3 I2 Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 VDD Z_neg ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 ZN Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   XNOR3_X4.                                                        *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:08 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT XNOR3_X4 A1 A2 A3 ZN VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VNW:P VPW:P VSS:G 
*.EQN ZN=!(!((!((A1 * A2) + !(A1 + A2)) * A3) + !(!((A1 * A2) + !(A1 + A2)) + A3)))
M_i_14 I A2 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_15 VSS A1 I VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 I2 I VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_0 net_0 A1 I2 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_1 VSS A2 net_0 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_18 I3 I2 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_19 VSS A3 I3 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_10 Z_neg I3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_8 net_2 A3 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_9 VSS I2 net_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_3 VSS Z_neg ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_2 ZN Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_1 VSS Z_neg ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_0 ZN Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_16 net_4 A2 I VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_17 VDD A1 net_4 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_5 net_1 I VDD VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_3 I2 A1 net_1 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_4 net_1 A2 I2 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_20 net_5 I2 I3 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_21 VDD A3 net_5 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_13 net_3 I3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11 Z_neg A3 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_12 net_3 I2 Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_3 VDD Z_neg ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_2 ZN Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 VDD Z_neg ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 ZN Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   XOR2_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:22 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT XOR2_X1 A1 A2 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=!((A1 * A2) + !(A1 + A2))
M_i_6 I A2 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_7 VSS A1 I VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_2 Z I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0 net_0 A1 Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1 VSS A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_8 net_2 A2 I VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_9 VDD A1 net_2 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_5 net_1 I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3 Z A1 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4 net_1 A2 Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   XOR2_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:24 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT XOR2_X2 A1 A2 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=!((A1 * A2) + !(A1 + A2))
M_i_8 net_2 A2 I VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_9 VSS A1 net_2 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_4 net_0 I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2 Z_neg A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 net_0 A2 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_10 I A2 VDD VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_11 VDD A1 I VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_7 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5 net_1 A1 Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 VDD A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   XOR2_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:24 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT XOR2_X4 A1 A2 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=!((A1 * A2) + !(A1 + A2))
M_i_8 net_2 A2 I VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_9 VSS A1 net_2 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_4 net_0 I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2 Z_neg A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 net_0 A2 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_10 I A2 VDD VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_11 VDD A1 I VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_7 Z_neg I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5 net_1 A1 Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 VDD A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_2 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   XOR3_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:05 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT XOR3_X1 A1 A2 A3 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=!((!((A1 * A2) + !(A1 + A2)) * A3) + !(!((A1 * A2) + !(A1 + A2)) + A3))
M_i_12 I A2 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_13 VSS A1 I VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 I2 I VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_0 net_0 A1 I2 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_1 VSS A2 net_0 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_16 I3 I2 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_17 VSS A3 I3 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_8 Z I3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6 net_2 A3 Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_7 VSS I2 net_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_14 net_4 A2 I VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_15 VDD A1 net_4 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_5 net_1 I VDD VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_3 I2 A1 net_1 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_4 net_1 A2 I2 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_18 net_5 I2 I3 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_19 VDD A3 net_5 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_11 net_3 I3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9 Z A3 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10 net_3 I2 Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   XOR3_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:07 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT XOR3_X2 A1 A2 A3 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=!((!((A1 * A2) + !(A1 + A2)) * A3) + !(!((A1 * A2) + !(A1 + A2)) + A3))
M_i_14 I A2 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_15 VSS A1 I VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 I2 I VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_0 net_0 A1 I2 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_1 VSS A2 net_0 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_18 net_5 I2 I3 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_19 VSS A3 net_5 VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_10 net_2 I3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_8 Z_neg A3 net_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_9 net_2 I2 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_1 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_16 net_4 A2 I VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_17 VDD A1 net_4 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_5 net_1 I VDD VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_3 I2 A1 net_1 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_4 net_1 A2 I2 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_20 I3 I2 VDD VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_21 VDD A3 I3 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_13 Z_neg I3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11 net_3 A3 Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_12 VDD I2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   XOR3_X4.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtcs026             *
* at 11:48:08 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT XOR3_X4 A1 A2 A3 Z VDD VNW VPW VSS 
*.PININFO A1:I A2:I A3:I Z:O VDD:P VNW:P VPW:P VSS:G 
*.EQN Z=!((!((A1 * A2) + !(A1 + A2)) * A3) + !(!((A1 * A2) + !(A1 + A2)) + A3))
M_i_14 I A2 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_15 VSS A1 I VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 I2 I VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_0 net_0 A1 I2 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_1 VSS A2 net_0 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_18 net_5 I2 I3 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_19 VSS A3 net_5 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_10 net_2 I3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_8 Z_neg A3 net_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_9 net_2 I2 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_3 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_2 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_1 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_16 net_4 A2 I VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_17 VDD A1 net_4 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_5 net_1 I VDD VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_3 I2 A1 net_1 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_4 net_1 A2 I2 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_20 I3 I2 VDD VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_21 VDD A3 I3 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_13 Z_neg I3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11 net_3 A3 Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_12 VDD I2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_3 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_2 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   ANTENNA.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Nanspice.                                                        *
*                                                                              *
* Written on scgtcs008             *
* at 16:34:20 on Tue, 18 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT ANTENNA I VDD VNW VPW VSS 
d0 VPW I np_6p0 0.2034p 1.85u $m=1
d1 I VNW pn_6p0 0.2034p 1.85u $m=1
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   ENDCAP.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* at 17:48:18 on Wed, 12 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT ENDCAP VDD VNW VPW VSS 
*.PININFO VDD:P VNW:P VPW:P VSS:G 

.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FILL_X1.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtgar01             *
* at 11:26:55 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT FILL_X1 VDD VNW VPW VSS 
*.PININFO VDD:P VNW:P VPW:P VSS:G 
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FILL_X2.                                                         *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtgar01             *
* at 11:26:55 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT FILL_X2 VDD VNW VPW VSS 
*.PININFO VDD:P VNW:P VPW:P VSS:G 
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FILL_X4.                                                           *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtgar01             *
* at 11:26:55 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT FILL_X4 VDD VNW VPW VSS 
*.PININFO VDD:P VNW:P VPW:P VSS:G 
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
*                                                                              *
* Cellname:   FILL_X8.                                                           *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtgar01             *
* at 11:26:55 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT FILL_X8 VDD VNW VPW VSS 
*.PININFO VDD:P VNW:P VPW:P VSS:G 
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FILL_X16.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtgar01             *
* at 11:26:55 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT FILL_X16 VDD VNW VPW VSS 
*.PININFO VDD:P VNW:P VPW:P VSS:G 
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FILL_X32.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtgar01             *
* at 11:26:55 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT FILL_X32 VDD VNW VPW VSS 
*.PININFO VDD:P VNW:P VPW:P VSS:G 
.ENDS 

********************************************************************************
*                                                                              *
* Cellname:   FILL_X64.                                                          *
*                                                                              *
* Technology: gf018.                                                           *
* Format:     Cdl.                                                             *
*                                                                              *
* Written on scgtgar01             *
* at 11:26:55 on Wed, 19 Mar 2014.                                             *
*                                                                              *
********************************************************************************
.SUBCKT FILL_X64 VDD VNW VPW VSS 
*.PININFO VDD:P VNW:P VPW:P VSS:G 
.ENDS 

********************************************************************************
*
* END
*
********************************************************************************
