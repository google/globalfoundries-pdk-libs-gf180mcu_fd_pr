************************************************************************
* auCdl Netlist:
* 
* Library Name:  TCG_Library
* Top Cell Name: diode_pw2dw_03v3
* View Name:     schematic
* Netlisted on:  Nov 24 09:06:01 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL vdd!

*.PIN vdd!

************************************************************************
* Library Name: TCG_Library
* Cell Name:    diode_pw2dw_03v3
* View Name:    schematic
************************************************************************

.SUBCKT diode_pw2dw_03v3 I1_0_0_0_0_0_R0_POS I1_0_1_0_0_0_R0_POS I1_0_2_0_0_0_R0_POS 
+ I1_1_0_0_0_0_R0_POS I1_1_1_0_0_0_R0_POS I1_1_2_0_0_0_R0_POS 
+ I1_2_0_0_0_0_R0_POS I1_2_1_0_0_0_R0_POS I1_2_2_0_0_0_R0_POS I1_default_POS 
+ vdd!
*.PININFO I1_0_0_0_0_0_R0_POS:I I1_0_1_0_0_0_R0_POS:I I1_0_2_0_0_0_R0_POS:I 
*.PININFO I1_1_0_0_0_0_R0_POS:I I1_1_1_0_0_0_R0_POS:I I1_1_2_0_0_0_R0_POS:I 
*.PININFO I1_2_0_0_0_0_R0_POS:I I1_2_1_0_0_0_R0_POS:I I1_2_2_0_0_0_R0_POS:I 
*.PININFO I1_default_POS:I vdd!:I
DI1_2_2_0_0_0_R0 I1_2_2_0_0_0_R0_POS vdd! diode_pw2dw_03v3 AREA=10n      PJ=400e-6    m=1
DI1_2_1_0_0_0_R0 I1_2_1_0_0_0_R0_POS vdd! diode_pw2dw_03v3 AREA=1.023n   PJ=220.46e-6 m=1
DI1_2_0_0_0_0_R0 I1_2_0_0_0_0_R0_POS vdd! diode_pw2dw_03v3 AREA=60p      PJ=201.2e-6  m=1
DI1_1_2_0_0_0_R0 I1_1_2_0_0_0_R0_POS vdd! diode_pw2dw_03v3 AREA=1.023n   PJ=220.46e-6 m=1
DI1_1_1_0_0_0_R0 I1_1_1_0_0_0_R0_POS vdd! diode_pw2dw_03v3 AREA=104.653p PJ=40.92e-6  m=1
DI1_1_0_0_0_0_R0 I1_1_0_0_0_0_R0_POS vdd! diode_pw2dw_03v3 AREA=6.138p   PJ=21.66e-6  m=1
DI1_0_2_0_0_0_R0 I1_0_2_0_0_0_R0_POS vdd! diode_pw2dw_03v3 AREA=60p      PJ=201.2e-6  m=1
DI1_0_1_0_0_0_R0 I1_0_1_0_0_0_R0_POS vdd! diode_pw2dw_03v3 AREA=6.138p   PJ=21.66e-6  m=1
DI1_0_0_0_0_0_R0 I1_0_0_0_0_0_R0_POS vdd! diode_pw2dw_03v3 AREA=627f     PJ=3.29e-6   m=1
DI1_default I1_default_POS vdd! diode_pw2dw_03v3 AREA=100e-12 PJ=40e-6 m=1
.ENDS

