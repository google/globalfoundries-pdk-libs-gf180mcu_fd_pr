* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

** Circuit sample_nfet_03v3

.subckt sample_nfet_03v3 I1_default_D I1_default_G I1_default_S vdd!
MI1_default I1_default_D I1_default_G I1_default_S vdd! nfet_03v3 m=1 w=360e-9
+ l=280n nf=1 as=158.4e-15 ad=158.4e-15 ps=1.6e-6 pd=1.6e-6 nrd=1.222222
+ nrs=1.222222 sa=0.440u sb=0.440u sd=0u dtemp=0 par=1
.ends

.end
