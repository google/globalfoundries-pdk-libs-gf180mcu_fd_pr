***************************
** CV netlist generation **
***************************
* Copyright 2022 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
Vb b 0 dc -3.0

.temp {{temp}}
.options tnom={{temp}}
      

xq1 0 b 0 0 {{device}}


.DC Vb 0 -3.0 -0.1

.control

save all @q.xq1.q0[cmu]
run 
print  @q.xq1.q0[cmu]

wrdata {{dirpath}}/cj_simulated/simulated_{{device}}_t{{temp}}_{{cap}}_{{corner}}.csv @q.xq1.q0[cmu]*1.0e15

.endc

** library calling

.include "../../../design.ngspice"
.lib "../../../sm141064.ngspice" bjt_{{corner}}


.end
