
*****************
** main netlist
*****************

Vcp c 0 dc 3
Vbp b 0 dc 1.2

xq1 c b 0 0 vnpn_10x10


*****************
** Analysis
*****************
.DC Vbp 0.2 1.2 0.01 Vcp 1 3 1
.STEP TEMP 25 -60 200
.print DC FORMAT=CSV file=result0.csv Vbp
.print DC FORMAT=CSV file=result0.csv {-I(Vbp)}
.print DC FORMAT=CSV file=result1.csv Vbp
.print DC FORMAT=CSV file=result1.csv {-I(Vcp)}

.include "../../../../design.xyce"
.lib "../../../../sm141064.xyce" bjt_typical

.end
