**************************
** res
**************************
* Copyright 2022 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

Vin top GND {{voltage}}
XR1 top {{terminals}} {{device}} r_width={{width}}u r_length={{length}}u m=1

.OP
.STEP TEMP 25 -60 200
.print DC {(V(top)*{{length}}u)/(-I(Vin)*{{width}}u)}


** library calling

.include "../../../design.xyce"
.lib "../../../sm141064.xyce" res_{{corner}}

.GLOBAL GND
.end
