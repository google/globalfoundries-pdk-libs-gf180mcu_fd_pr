.SUBCKT gf180mcu_fd_io__bi_24t A CS DVDD DVSS IE OE PAD PD PU SL VDD VSS Y
R0 n9 VDD $SUB=VDD $[ppolyf_u] $W=800e-9 $L=1.6e-6 m=1.0 r=907.859 par=1
R1 n11 VDD $SUB=VDD $[ppolyf_u] $W=800e-9 $L=1.6e-6 m=1.0 r=907.859 par=1
C2 DVDD DVSS $[cap_nmos_06v0] m=4.0 l=3e-6 w=3e-6
C3 DVDD DVSS $[cap_nmos_06v0] m=8.0 l=1.5e-6 w=5e-6
M4 n43 n32 DVSS DVSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 ad=780e-15 
+ ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9 
+ sd=520e-9 dtemp=0.0 par=1
M5 n56 IE VSS VSS nfet_06v0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 ad=660e-15 
+ ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M6 n32 n56 DVSS DVSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 ad=780e-15 
+ ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9 
+ sd=520e-9 dtemp=0.0 par=1
M7 n43 n32 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 ad=1.56e-12 
+ ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 sb=440e-9 
+ sd=520e-9 dtemp=0.0 par=1
M8 n56 IE VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 ad=1.32e-12 
+ ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M9 n32 n56 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 ad=1.56e-12 
+ ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 sb=440e-9 
+ sd=520e-9 dtemp=0.0 par=1
M10 n49 n33 DVSS DVSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 ad=780e-15 
+ ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9 
+ sd=520e-9 dtemp=0.0 par=1
M11 n64 CS VSS VSS nfet_06v0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M12 n33 n64 DVSS DVSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 ad=780e-15 
+ ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9 
+ sd=520e-9 dtemp=0.0 par=1
M13 n49 n33 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M14 n64 CS VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M15 n33 n64 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M16 n47 n35 DVSS DVSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 ad=780e-15 
+ ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9 
+ sd=520e-9 dtemp=0.0 par=1
M17 n72 n36 VSS VSS nfet_06v0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M18 n35 n72 DVSS DVSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 ad=780e-15 
+ ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9 
+ sd=520e-9 dtemp=0.0 par=1
M19 n47 n35 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M20 n72 n36 VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M21 n35 n72 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M22 n51 n38 DVSS DVSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 ad=780e-15 
+ ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9 
+ sd=520e-9 dtemp=0.0 par=1
M23 n80 n34 VSS VSS nfet_06v0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M24 n38 n80 DVSS DVSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 ad=780e-15 
+ ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9 
+ sd=520e-9 dtemp=0.0 par=1
M25 n51 n38 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M26 n80 n34 VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M27 n38 n80 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
D28 PD VDD diode_pd2nw_06v0 m=1.0 AREA=1e-12 PJ=4e-6
D29 IE VDD diode_pd2nw_06v0 m=1.0 AREA=1e-12 PJ=4e-6
D30 CS VDD diode_pd2nw_06v0 m=1.0 AREA=1e-12 PJ=4e-6
D31 PU VDD diode_pd2nw_06v0 m=1.0 AREA=1e-12 PJ=4e-6
M32 n88 n33 DVDD DVDD pfet_06v0 m=1.0 w=8e-6 l=700e-9 nf=1.0 as=3.52e-12 
+ ad=3.52e-12 ps=16.88e-6 pd=16.88e-6 nrd=55e-3 nrs=55e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M33 DVDD n33 n89 DVDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M34 n90 n21 DVDD DVDD pfet_06v0 m=1.0 w=3.8e-6 l=700e-9 nf=1.0 as=1.672e-12 
+ ad=1.672e-12 ps=8.48e-6 pd=8.48e-6 nrd=115.789e-3 nrs=115.789e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M35 DVSS n89 n90 DVDD pfet_06v0 m=1.0 w=3.8e-6 l=700e-9 nf=1.0 as=1.672e-12 
+ ad=1.672e-12 ps=8.48e-6 pd=8.48e-6 nrd=115.789e-3 nrs=115.789e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M36 n50 n32 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M37 n50 n88 n85 DVDD pfet_06v0 m=1.0 w=2e-6 l=700e-9 nf=1.0 as=880e-15 ad=880e-15 
+ ps=4.88e-6 pd=4.88e-6 nrd=220e-3 nrs=220e-3 sa=440e-9 sb=440e-9 sd=0.0 
+ dtemp=0.0 par=1
M38 n50 n88 n89 DVDD pfet_06v0 m=1.0 w=2e-6 l=700e-9 nf=1.0 as=880e-15 ad=880e-15 
+ ps=4.88e-6 pd=4.88e-6 nrd=220e-3 nrs=220e-3 sa=440e-9 sb=440e-9 sd=0.0 
+ dtemp=0.0 par=1
M39 n50 n21 n90 DVDD pfet_06v0 m=1.0 w=4.3e-6 l=700e-9 nf=1.0 as=1.892e-12 
+ ad=1.892e-12 ps=9.48e-6 pd=9.48e-6 nrd=102.326e-3 nrs=102.326e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M40 n95 n32 DVSS DVSS nfet_06v0 m=1.0 w=16e-6 l=700e-9 nf=1.0 as=7.04e-12 
+ ad=7.04e-12 ps=32.88e-6 pd=32.88e-6 nrd=27.5e-3 nrs=27.5e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M41 n87 n21 n95 DVSS nfet_06v0 m=1.0 w=10.6e-6 l=700e-9 nf=1.0 as=4.664e-12 
+ ad=4.664e-12 ps=22.08e-6 pd=22.08e-6 nrd=41.509e-3 nrs=41.509e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M42 n50 n21 n87 DVSS nfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M43 n88 n33 DVSS DVSS nfet_06v0 m=1.0 w=4e-6 l=700e-9 nf=1.0 as=1.76e-12 
+ ad=1.76e-12 ps=8.88e-6 pd=8.88e-6 nrd=110e-3 nrs=110e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M44 n50 n33 n85 DVSS nfet_06v0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M45 n50 n33 n89 DVSS nfet_06v0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M46 DVDD n85 n87 DVSS nfet_06v0 m=1.0 w=1.3e-6 l=700e-9 nf=1.0 as=572e-15 
+ ad=572e-15 ps=3.48e-6 pd=3.48e-6 nrd=338.462e-3 nrs=338.462e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M47 DVSS n88 n85 DVSS nfet_06v0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M48 n103 n50 DVDD DVDD pfet_06v0 m=1.0 w=2e-6 l=700e-9 nf=1.0 as=880e-15 ad=880e-15 
+ ps=4.88e-6 pd=4.88e-6 nrd=220e-3 nrs=220e-3 sa=440e-9 sb=440e-9 sd=0.0 
+ dtemp=0.0 par=1
M49 n100 n103 VDD VDD pfet_06v0 m=1.0 w=10e-6 l=700e-9 nf=1.0 as=4.4e-12 
+ ad=4.4e-12 ps=20.88e-6 pd=20.88e-6 nrd=44e-3 nrs=44e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M50 Y n100 VDD VDD pfet_06v0 m=1.0 w=21e-6 l=700e-9 nf=1.0 as=9.24e-12 
+ ad=9.24e-12 ps=42.88e-6 pd=42.88e-6 nrd=20.952e-3 nrs=20.952e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M51 n103 n50 DVSS DVSS nfet_06v0 m=1.0 w=8e-6 l=700e-9 nf=1.0 as=3.52e-12 
+ ad=3.52e-12 ps=16.88e-6 pd=16.88e-6 nrd=55e-3 nrs=55e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M52 Y n100 VSS VSS nfet_06v0 m=1.0 w=9e-6 l=700e-9 nf=1.0 as=3.96e-12 
+ ad=3.96e-12 ps=18.88e-6 pd=18.88e-6 nrd=48.889e-3 nrs=48.889e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M53 n100 n103 VSS VSS nfet_06v0 m=1.0 w=2.5e-6 l=700e-9 nf=1.0 as=1.1e-12 
+ ad=1.1e-12 ps=5.88e-6 pd=5.88e-6 nrd=176e-3 nrs=176e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M54 n36 n110 VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M55 n36 PU VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 ad=1.32e-12 
+ ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M56 n111 PU VSS VSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M57 n36 n110 n111 VSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M58 n34 PD VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 ad=1.32e-12 
+ ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 sb=440e-9 
+ sd=0.0 dtemp=0.0 par=1
M59 n34 n110 VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M60 n117 n110 VSS VSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M61 n34 PD n117 VSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M62 n123 n129 n110 VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M63 PU PD n110 VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M64 n129 PD VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M65 n123 PU VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M66 n123 PD n110 VSS nfet_06v0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M67 PU n129 n110 VSS nfet_06v0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M68 n129 PD VSS VSS nfet_06v0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M69 n123 PU VSS VSS nfet_06v0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
R70 n21 n132 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=23e-6 m=1.0 r=9.94533e3 par=1
R71 n132 n131 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
R72 n131 n130 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
R73 n130 n133 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
R74 n133 n138 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
R75 n138 n137 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
R76 n137 n134 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
R77 n134 n135 $SUB=DVDD $[ppolyf_u] $W=800e-9 $L=35.7e-6 m=1.0 r=15.3065e3 par=1
M78 n135 n51 DVSS DVSS nfet_06v0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M79 n135 n35 DVDD DVDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
D80 DVSS n21 diode_nd2ps_06v0 m=2.0 AREA=20e-12 PJ=42e-6
D81 n21 DVDD diode_pd2nw_06v0 m=2.0 AREA=20e-12 PJ=42e-6
R82 PAD n21 $SUB=DVDD $[ppolyf_u] $W=2.5e-6 $L=2.8e-6 m=1.0 r=432.59 par=1
R83 PAD n21 $SUB=DVDD $[ppolyf_u] $W=2.5e-6 $L=2.8e-6 m=1.0 r=449.157 par=1
R84 PAD n21 $SUB=DVDD $[ppolyf_u] $W=2.5e-6 $L=2.8e-6 m=1.0 r=432.59 par=1
R85 PAD n21 $SUB=DVDD $[ppolyf_u] $W=2.5e-6 $L=2.8e-6 m=1.0 r=449.157 par=1
M86 n183 n191 DVSS DVSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M87 n153 n183 DVSS DVSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M88 n188 OE VSS VSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M89 n191 A n188 VSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M90 n183 n191 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M91 n153 n183 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M92 n191 OE VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M93 n191 A VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M94 PAD n157 DVDD DVDD pfet_06v0_dss m=1.0 w=120e-6 l=700e-9 nf=2.0 s_sab=280e-9 
+ d_sab=2.78e-6 par=1 dtemp=0.0
M95 PAD n165 DVDD DVDD pfet_06v0_dss m=1.0 w=60e-6 l=700e-9 nf=1.0 s_sab=280e-9 
+ d_sab=2.78e-6 par=1 dtemp=0.0
M96 PAD n172 DVSS DVSS nfet_06v0_dss m=1.0 w=37e-6 l=800e-9 nf=1.0 s_sab=280e-9 
+ d_sab=3.78e-6 par=1 dtemp=0.0
M97 PAD n169 DVSS DVSS nfet_06v0_dss m=1.0 w=37e-6 l=800e-9 nf=1.0 s_sab=280e-9 
+ d_sab=3.78e-6 par=1 dtemp=0.0
M98 PAD n158 DVDD DVDD pfet_06v0_dss m=1.0 w=120e-6 l=700e-9 nf=2.0 s_sab=280e-9 
+ d_sab=2.78e-6 par=1 dtemp=0.0
M99 PAD n164 DVDD DVDD pfet_06v0_dss m=1.0 w=60e-6 l=700e-9 nf=1.0 s_sab=280e-9 
+ d_sab=2.78e-6 par=1 dtemp=0.0
M100 PAD n173 DVSS DVSS nfet_06v0_dss m=1.0 w=37e-6 l=800e-9 nf=1.0 s_sab=280e-9 
+ d_sab=3.78e-6 par=1 dtemp=0.0
M101 PAD n168 DVSS DVSS nfet_06v0_dss m=1.0 w=37e-6 l=800e-9 nf=1.0 s_sab=280e-9 
+ d_sab=3.78e-6 par=1 dtemp=0.0
M102 PAD n161 DVDD DVDD pfet_06v0_dss m=1.0 w=120e-6 l=700e-9 nf=2.0 s_sab=280e-9 
+ d_sab=2.78e-6 par=1 dtemp=0.0
M103 PAD n166 DVDD DVDD pfet_06v0_dss m=1.0 w=60e-6 l=700e-9 nf=1.0 s_sab=280e-9 
+ d_sab=2.78e-6 par=1 dtemp=0.0
M104 PAD n171 DVSS DVSS nfet_06v0_dss m=1.0 w=37e-6 l=800e-9 nf=1.0 s_sab=280e-9 
+ d_sab=3.78e-6 par=1 dtemp=0.0
M105 PAD n170 DVSS DVSS nfet_06v0_dss m=1.0 w=37e-6 l=800e-9 nf=1.0 s_sab=280e-9 
+ d_sab=3.78e-6 par=1 dtemp=0.0
M106 PAD n162 DVDD DVDD pfet_06v0_dss m=1.0 w=120e-6 l=700e-9 nf=2.0 s_sab=280e-9 
+ d_sab=2.78e-6 par=1 dtemp=0.0
M107 PAD n163 DVDD DVDD pfet_06v0_dss m=1.0 w=60e-6 l=700e-9 nf=1.0 s_sab=280e-9 
+ d_sab=2.78e-6 par=1 dtemp=0.0
M108 PAD n174 DVSS DVSS nfet_06v0_dss m=1.0 w=37e-6 l=800e-9 nf=1.0 s_sab=280e-9 
+ d_sab=3.78e-6 par=1 dtemp=0.0
M109 PAD n167 DVSS DVSS nfet_06v0_dss m=1.0 w=37e-6 l=800e-9 nf=1.0 s_sab=280e-9 
+ d_sab=3.78e-6 par=1 dtemp=0.0
D110 A VDD diode_pd2nw_06v0 m=1.0 AREA=1e-12 PJ=4e-6
D111 SL VDD diode_pd2nw_06v0 m=1.0 AREA=1e-12 PJ=4e-6
M112 n159 n160 DVSS DVSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M113 n291 SL VSS VSS nfet_06v0 m=1.0 w=1.5e-6 l=700e-9 nf=1.0 as=660e-15 
+ ad=660e-15 ps=3.88e-6 pd=3.88e-6 nrd=293.333e-3 nrs=293.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M114 n160 n291 DVSS DVSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=2.0 as=1.32e-12 
+ ad=780e-15 ps=7.76e-6 pd=4.04e-6 nrd=86.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M115 n159 n160 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
M116 n291 SL VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M117 n160 n291 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=2.0 as=2.64e-12 
+ ad=1.56e-12 ps=13.76e-6 pd=7.04e-6 nrd=43.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=520e-9 dtemp=0.0 par=1
D118 VSS n9 diode_pd2nw_06v0 m=1.0 AREA=230.4e-15 PJ=1.92e-6
D119 VSS OE diode_pd2nw_06v0 m=1.0 AREA=230.4e-15 PJ=1.92e-6
M120 n304 n9 VSS VSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M121 n295 OE n304 VSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M122 n156 n152 DVSS DVSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M123 n152 n295 DVSS DVSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M124 n295 n9 VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M125 n295 OE VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M126 n156 n152 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M127 n152 n295 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
D128 VSS n11 diode_pd2nw_06v0 m=1.0 AREA=230.4e-15 PJ=1.92e-6
D129 VSS OE diode_pd2nw_06v0 m=1.0 AREA=230.4e-15 PJ=1.92e-6
M130 n314 n11 VSS VSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M131 n305 OE n314 VSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M132 n151 n150 DVSS DVSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M133 n150 n305 DVSS DVSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M134 n305 n11 VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M135 n305 OE VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M136 n151 n150 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M137 n150 n305 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
D138 VSS VDD diode_pd2nw_06v0 m=1.0 AREA=230.4e-15 PJ=1.92e-6
D139 VSS OE diode_pd2nw_06v0 m=1.0 AREA=230.4e-15 PJ=1.92e-6
M140 n324 VDD VSS VSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M141 n315 OE n324 VSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M142 n148 n147 DVSS DVSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M143 n147 n315 DVSS DVSS nfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M144 n315 VDD VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M145 n315 OE VDD VDD pfet_06v0 m=1.0 w=3e-6 l=700e-9 nf=1.0 as=1.32e-12 
+ ad=1.32e-12 ps=6.88e-6 pd=6.88e-6 nrd=146.667e-3 nrs=146.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M146 n148 n147 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M147 n147 n315 DVDD DVDD pfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M148 n163 n159 n162 DVSS nfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M149 n162 DVDD n163 DVSS nfet_06v0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15 
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M150 n167 n325 DVSS DVSS nfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M151 n174 n325 DVSS DVSS nfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M152 n163 n330 DVSS DVSS nfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M153 n330 n153 DVSS DVSS nfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M154 n330 n156 DVSS DVSS nfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M155 n325 n152 n330 DVSS nfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M156 n167 n160 n174 DVDD pfet_06v0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M157 n325 n152 DVDD DVDD pfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M158 n163 n330 DVDD DVDD pfet_06v0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M159 n174 n325 DVDD DVDD pfet_06v0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M160 n167 DVSS n174 DVDD pfet_06v0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15 
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M161 n325 n153 DVDD DVDD pfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M162 n330 n156 n325 DVDD pfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M163 n162 n330 DVDD DVDD pfet_06v0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M164 n164 n159 n158 DVSS nfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M165 n158 DVDD n164 DVSS nfet_06v0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15 
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M166 n168 n338 DVSS DVSS nfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M167 n173 n338 DVSS DVSS nfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M168 n164 n343 DVSS DVSS nfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M169 n343 n153 DVSS DVSS nfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M170 n343 n151 DVSS DVSS nfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M171 n338 n150 n343 DVSS nfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M172 n168 n160 n173 DVDD pfet_06v0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M173 n338 n150 DVDD DVDD pfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M174 n164 n343 DVDD DVDD pfet_06v0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M175 n173 n338 DVDD DVDD pfet_06v0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M176 n168 DVSS n173 DVDD pfet_06v0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15 
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M177 n338 n153 DVDD DVDD pfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M178 n343 n151 n338 DVDD pfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M179 n158 n343 DVDD DVDD pfet_06v0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M180 n165 n159 n157 DVSS nfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M181 n157 DVDD n165 DVSS nfet_06v0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15 
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M182 n169 n351 DVSS DVSS nfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M183 n172 n351 DVSS DVSS nfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M184 n165 n356 DVSS DVSS nfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M185 n356 n153 DVSS DVSS nfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M186 n356 n151 DVSS DVSS nfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M187 n351 n150 n356 DVSS nfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M188 n169 n160 n172 DVDD pfet_06v0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M189 n351 n150 DVDD DVDD pfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M190 n165 n356 DVDD DVDD pfet_06v0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M191 n172 n351 DVDD DVDD pfet_06v0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M192 n169 DVSS n172 DVDD pfet_06v0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15 
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M193 n351 n153 DVDD DVDD pfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M194 n356 n151 n351 DVDD pfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M195 n157 n356 DVDD DVDD pfet_06v0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M196 n166 n159 n161 DVSS nfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M197 n161 DVDD n166 DVSS nfet_06v0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15 
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M198 n170 n364 DVSS DVSS nfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M199 n171 n364 DVSS DVSS nfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M200 n166 n369 DVSS DVSS nfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M201 n369 n153 DVSS DVSS nfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M202 n369 n148 DVSS DVSS nfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M203 n364 n147 n369 DVSS nfet_06v0 m=1.0 w=6e-6 l=700e-9 nf=1.0 as=2.64e-12 
+ ad=2.64e-12 ps=12.88e-6 pd=12.88e-6 nrd=73.333e-3 nrs=73.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M204 n170 n160 n171 DVDD pfet_06v0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M205 n364 n147 DVDD DVDD pfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M206 n166 n369 DVDD DVDD pfet_06v0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M207 n171 n364 DVDD DVDD pfet_06v0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M208 n170 DVSS n171 DVDD pfet_06v0 m=1.0 w=1.2e-6 l=700e-9 nf=1.0 as=528e-15 
+ ad=528e-15 ps=3.28e-6 pd=3.28e-6 nrd=366.667e-3 nrs=366.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M209 n364 n153 DVDD DVDD pfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M210 n369 n148 n364 DVDD pfet_06v0 m=1.0 w=12e-6 l=700e-9 nf=1.0 as=5.28e-12 
+ ad=5.28e-12 ps=24.88e-6 pd=24.88e-6 nrd=36.667e-3 nrs=36.667e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
M211 n161 n369 DVDD DVDD pfet_06v0 m=1.0 w=24e-6 l=700e-9 nf=1.0 as=10.56e-12 
+ ad=10.56e-12 ps=48.88e-6 pd=48.88e-6 nrd=18.333e-3 nrs=18.333e-3 sa=440e-9 
+ sb=440e-9 sd=0.0 dtemp=0.0 par=1
.ENDS
