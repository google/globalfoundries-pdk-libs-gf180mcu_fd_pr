************************************************************************
* auCdl Netlist:
* 
* Library Name:  TCG_library_2
* Top Cell Name: sample_gppmos_6p0_dw_sab
* View Name:     schematic
* Netlisted on:  Sep 10 16:24:13 2021
************************************************************************

*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL sub!

*.PIN sub!

************************************************************************
* Library Name: TCG_library_2
* Cell Name:    sample_gppmos_6p0_dw_sab
* View Name:    schematic
************************************************************************

.SUBCKT sample_gppmos_6p0_dw_sab I1_default_D I1_lin_default_d_sab_0_R0_D 
+ I1_lin_default_d_sab_1_R0_D I1_lin_default_d_sab_2_R0_D 
+ I1_lin_default_d_sab_3_R0_D I1_lin_default_d_sab_4_R0_D 
+ I1_lin_default_d_sab_5_R0_D I1_lin_default_d_sab_6_R0_D 
+ I1_lin_default_d_sab_7_R0_D I1_lin_default_d_sab_8_R0_D 
+ I1_lin_default_d_sab_9_R0_D I1_lin_default_gns_0_R0_D 
+ I1_lin_default_gns_1_R0_D I1_lin_default_guardRing_0_R0_D 
+ I1_lin_default_l_0_R0_D I1_lin_default_l_1_R0_D I1_lin_default_l_2_R0_D 
+ I1_lin_default_l_3_R0_D I1_lin_default_l_4_R0_D I1_lin_default_l_5_R0_D 
+ I1_lin_default_l_6_R0_D I1_lin_default_l_7_R0_D I1_lin_default_l_8_R0_D 
+ I1_lin_default_l_9_R0_D I1_lin_default_l_10_R0_D I1_lin_default_l_11_R0_D 
+ I1_lin_default_l_12_R0_D I1_lin_default_l_13_R0_D I1_lin_default_l_14_R0_D 
+ I1_lin_default_l_15_R0_D I1_lin_default_m_0_R0_D I1_lin_default_m_1_R0_D 
+ I1_lin_default_m_2_R0_D I1_lin_default_nf_0_R0_D I1_lin_default_nf_1_R0_D 
+ I1_lin_default_nf_2_R0_D I1_lin_default_nf_3_R0_D I1_lin_default_nf_4_R0_D 
+ I1_lin_default_nf_5_R0_D I1_lin_default_nf_6_R0_D 
+ I1_lin_default_psub_tap_0_R0_D I1_lin_default_s_sab_0_R0_D 
+ I1_lin_default_s_sab_1_R0_D I1_lin_default_s_sab_2_R0_D 
+ I1_lin_default_s_sab_3_R0_D I1_lin_default_s_sab_4_R0_D 
+ I1_lin_default_s_sab_5_R0_D I1_lin_default_s_sab_6_R0_D 
+ I1_lin_default_s_sab_7_R0_D I1_lin_default_strapSD_0_R0_D 
+ I1_lin_default_wf_0_R0_D I1_lin_default_wf_1_R0_D I1_lin_default_wf_2_R0_D 
+ I1_lin_default_wf_3_R0_D I1_lin_default_wf_4_R0_D sub!
*.PININFO I1_default_D:I I1_lin_default_d_sab_0_R0_D:I 
*.PININFO I1_lin_default_d_sab_1_R0_D:I I1_lin_default_d_sab_2_R0_D:I 
*.PININFO I1_lin_default_d_sab_3_R0_D:I I1_lin_default_d_sab_4_R0_D:I 
*.PININFO I1_lin_default_d_sab_5_R0_D:I I1_lin_default_d_sab_6_R0_D:I 
*.PININFO I1_lin_default_d_sab_7_R0_D:I I1_lin_default_d_sab_8_R0_D:I 
*.PININFO I1_lin_default_d_sab_9_R0_D:I I1_lin_default_gns_0_R0_D:I 
*.PININFO I1_lin_default_gns_1_R0_D:I I1_lin_default_guardRing_0_R0_D:I 
*.PININFO I1_lin_default_l_0_R0_D:I I1_lin_default_l_1_R0_D:I 
*.PININFO I1_lin_default_l_2_R0_D:I I1_lin_default_l_3_R0_D:I 
*.PININFO I1_lin_default_l_4_R0_D:I I1_lin_default_l_5_R0_D:I 
*.PININFO I1_lin_default_l_6_R0_D:I I1_lin_default_l_7_R0_D:I 
*.PININFO I1_lin_default_l_8_R0_D:I I1_lin_default_l_9_R0_D:I 
*.PININFO I1_lin_default_l_10_R0_D:I I1_lin_default_l_11_R0_D:I 
*.PININFO I1_lin_default_l_12_R0_D:I I1_lin_default_l_13_R0_D:I 
*.PININFO I1_lin_default_l_14_R0_D:I I1_lin_default_l_15_R0_D:I 
*.PININFO I1_lin_default_m_0_R0_D:I I1_lin_default_m_1_R0_D:I 
*.PININFO I1_lin_default_m_2_R0_D:I I1_lin_default_nf_0_R0_D:I 
*.PININFO I1_lin_default_nf_1_R0_D:I I1_lin_default_nf_2_R0_D:I 
*.PININFO I1_lin_default_nf_3_R0_D:I I1_lin_default_nf_4_R0_D:I 
*.PININFO I1_lin_default_nf_5_R0_D:I I1_lin_default_nf_6_R0_D:I 
*.PININFO I1_lin_default_psub_tap_0_R0_D:I I1_lin_default_s_sab_0_R0_D:I 
*.PININFO I1_lin_default_s_sab_1_R0_D:I I1_lin_default_s_sab_2_R0_D:I 
*.PININFO I1_lin_default_s_sab_3_R0_D:I I1_lin_default_s_sab_4_R0_D:I 
*.PININFO I1_lin_default_s_sab_5_R0_D:I I1_lin_default_s_sab_6_R0_D:I 
*.PININFO I1_lin_default_s_sab_7_R0_D:I I1_lin_default_strapSD_0_R0_D:I 
*.PININFO I1_lin_default_wf_0_R0_D:I I1_lin_default_wf_1_R0_D:I 
*.PININFO I1_lin_default_wf_2_R0_D:I I1_lin_default_wf_3_R0_D:I 
*.PININFO I1_lin_default_wf_4_R0_D:I sub!:I
MI1_lin_default_wf_4_R0 I1_lin_default_wf_4_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=720.000u l=0.7u nf=18 s_sab=0.28u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_wf_3_R0 I1_lin_default_wf_3_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=622.080u l=0.7u nf=18 s_sab=0.28u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_wf_2_R0 I1_lin_default_wf_2_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=518.400u l=0.7u nf=18 s_sab=0.28u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_wf_1_R0 I1_lin_default_wf_1_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=432.000u l=0.7u nf=18 s_sab=0.28u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_wf_0_R0 I1_lin_default_wf_0_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=360.000u l=0.7u nf=18 s_sab=0.28u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_l_15_R0 I1_lin_default_l_15_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=10.000u nf=18 s_sab=0.28u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_l_14_R0 I1_lin_default_l_14_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=8.985u nf=18 s_sab=0.28u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_l_13_R0 I1_lin_default_l_13_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=7.490u nf=18 s_sab=0.28u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_l_12_R0 I1_lin_default_l_12_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=6.240u nf=18 s_sab=0.28u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_l_11_R0 I1_lin_default_l_11_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=5.200u nf=18 s_sab=0.28u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_l_10_R0 I1_lin_default_l_10_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=4.335u nf=18 s_sab=0.28u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_l_9_R0 I1_lin_default_l_9_R0_D sub! sub! sub! pmos_6p0_dw_sab 
+ m=1 w=450u l=3.610u nf=18 s_sab=0.28u d_sab=2.78u par=1 dtemp=0
MI1_lin_default_l_8_R0 I1_lin_default_l_8_R0_D sub! sub! sub! pmos_6p0_dw_sab 
+ m=1 w=450u l=3.010u nf=18 s_sab=0.28u d_sab=2.78u par=1 dtemp=0
MI1_lin_default_l_7_R0 I1_lin_default_l_7_R0_D sub! sub! sub! pmos_6p0_dw_sab 
+ m=1 w=450u l=2.510u nf=18 s_sab=0.28u d_sab=2.78u par=1 dtemp=0
MI1_lin_default_l_6_R0 I1_lin_default_l_6_R0_D sub! sub! sub! pmos_6p0_dw_sab 
+ m=1 w=450u l=2.090u nf=18 s_sab=0.28u d_sab=2.78u par=1 dtemp=0
MI1_lin_default_l_5_R0 I1_lin_default_l_5_R0_D sub! sub! sub! pmos_6p0_dw_sab 
+ m=1 w=450u l=1.740u nf=18 s_sab=0.28u d_sab=2.78u par=1 dtemp=0
MI1_lin_default_l_4_R0 I1_lin_default_l_4_R0_D sub! sub! sub! pmos_6p0_dw_sab 
+ m=1 w=450u l=1.450u nf=18 s_sab=0.28u d_sab=2.78u par=1 dtemp=0
MI1_lin_default_l_3_R0 I1_lin_default_l_3_R0_D sub! sub! sub! pmos_6p0_dw_sab 
+ m=1 w=450u l=1.210u nf=18 s_sab=0.28u d_sab=2.78u par=1 dtemp=0
MI1_lin_default_l_2_R0 I1_lin_default_l_2_R0_D sub! sub! sub! pmos_6p0_dw_sab 
+ m=1 w=450u l=1.010u nf=18 s_sab=0.28u d_sab=2.78u par=1 dtemp=0
MI1_lin_default_l_1_R0 I1_lin_default_l_1_R0_D sub! sub! sub! pmos_6p0_dw_sab 
+ m=1 w=450u l=0.840u nf=18 s_sab=0.28u d_sab=2.78u par=1 dtemp=0
MI1_lin_default_l_0_R0 I1_lin_default_l_0_R0_D sub! sub! sub! pmos_6p0_dw_sab 
+ m=1 w=450u l=0.700u nf=18 s_sab=0.28u d_sab=2.78u par=1 dtemp=0
MI1_lin_default_d_sab_9_R0 I1_lin_default_d_sab_9_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.28u d_sab=3.780u par=1 
+ dtemp=0
MI1_lin_default_d_sab_8_R0 I1_lin_default_d_sab_8_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.28u d_sab=3.355u par=1 
+ dtemp=0
MI1_lin_default_d_sab_7_R0 I1_lin_default_d_sab_7_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.28u d_sab=2.795u par=1 
+ dtemp=0
MI1_lin_default_d_sab_6_R0 I1_lin_default_d_sab_6_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.28u d_sab=2.330u par=1 
+ dtemp=0
MI1_lin_default_d_sab_5_R0 I1_lin_default_d_sab_5_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.28u d_sab=1.940u par=1 
+ dtemp=0
MI1_lin_default_d_sab_4_R0 I1_lin_default_d_sab_4_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.28u d_sab=1.615u par=1 
+ dtemp=0
MI1_lin_default_d_sab_3_R0 I1_lin_default_d_sab_3_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.28u d_sab=1.350u par=1 
+ dtemp=0
MI1_lin_default_d_sab_2_R0 I1_lin_default_d_sab_2_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.28u d_sab=1.125u par=1 
+ dtemp=0
MI1_lin_default_d_sab_1_R0 I1_lin_default_d_sab_1_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.28u d_sab=0.935u par=1 
+ dtemp=0
MI1_lin_default_d_sab_0_R0 I1_lin_default_d_sab_0_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.28u d_sab=0.780u par=1 
+ dtemp=0
MI1_lin_default_s_sab_7_R0 I1_lin_default_s_sab_7_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.780u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_s_sab_6_R0 I1_lin_default_s_sab_6_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.655u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_s_sab_5_R0 I1_lin_default_s_sab_5_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.545u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_s_sab_4_R0 I1_lin_default_s_sab_4_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.455u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_s_sab_3_R0 I1_lin_default_s_sab_3_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.380u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_s_sab_2_R0 I1_lin_default_s_sab_2_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.315u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_s_sab_1_R0 I1_lin_default_s_sab_1_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.265u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_s_sab_0_R0 I1_lin_default_s_sab_0_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.220u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_nf_6_R0 I1_lin_default_nf_6_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=600.000u l=0.7u nf=24 s_sab=0.28u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_nf_5_R0 I1_lin_default_nf_5_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=550.000u l=0.7u nf=22 s_sab=0.28u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_nf_4_R0 I1_lin_default_nf_4_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=500.000u l=0.7u nf=20 s_sab=0.28u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_nf_3_R0 I1_lin_default_nf_3_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450.000u l=0.7u nf=18 s_sab=0.28u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_nf_2_R0 I1_lin_default_nf_2_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=400.000u l=0.7u nf=16 s_sab=0.28u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_nf_1_R0 I1_lin_default_nf_1_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=350.000u l=0.7u nf=14 s_sab=0.28u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_nf_0_R0 I1_lin_default_nf_0_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=300.000u l=0.7u nf=12 s_sab=0.28u d_sab=2.78u par=1 
+ dtemp=0
MI1_lin_default_m_2_R0 I1_lin_default_m_2_R0_D sub! sub! sub! pmos_6p0_dw_sab 
+ m=3 w=450u l=0.7u nf=18 s_sab=0.28u d_sab=2.78u par=3 dtemp=0
MI1_lin_default_m_1_R0 I1_lin_default_m_1_R0_D sub! sub! sub! pmos_6p0_dw_sab 
+ m=2 w=450u l=0.7u nf=18 s_sab=0.28u d_sab=2.78u par=2 dtemp=0
MI1_lin_default_m_0_R0 I1_lin_default_m_0_R0_D sub! sub! sub! pmos_6p0_dw_sab 
+ m=1 w=450u l=0.7u nf=18 s_sab=0.28u d_sab=2.78u par=1 dtemp=0
MI1_lin_default_gns_1_R0 I1_lin_default_gns_1_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0 d_sab=2.78u par=1 dtemp=0
MI1_lin_default_gns_0_R0 I1_lin_default_gns_0_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.28u d_sab=2.78u par=1 dtemp=0
MI1_lin_default_guardRing_0_R0 I1_lin_default_guardRing_0_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.28u d_sab=2.78u par=1 dtemp=0
MI1_lin_default_strapSD_0_R0 I1_lin_default_strapSD_0_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.28u d_sab=2.78u par=1 dtemp=0
MI1_lin_default_psub_tap_0_R0 I1_lin_default_psub_tap_0_R0_D sub! sub! sub! 
+ pmos_6p0_dw_sab m=1 w=450u l=0.7u nf=18 s_sab=0.28u d_sab=2.78u par=1 dtemp=0
MI1_default I1_default_D sub! sub! sub! pmos_6p0_dw_sab m=1 w=450u l=0.7u 
+ nf=18 s_sab=0.28u d_sab=2.78u par=1 dtemp=0
.ENDS

