* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

**************************************
* Revision: 1.0
**************************************


*.SCALE METER

.SUBCKT power_route_04
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_PSUB_I01
** N=2765 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_PSUB_I06
** N=2653 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_PSUB$$47122476
** N=5 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nfet_05v0_I08
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pfet_05v0_I09 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 pfet_05v0 L=6e-07 W=6.81e-06 AD=2.9964e-12 AS=2.9964e-12 PD=1.45e-05 PS=1.45e-05 NRD=0.0646109 NRS=0.0646109 m=1 nf=1 $X=0 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT pmos_1p2$$46889004 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
X0 1 2 3 4 pfet_05v0_I09 $T=-155 0 0 0 $X=-1195 $Y=-620
.ENDS
***************************************
.SUBCKT nfet_05v0_I12 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 nfet_05v0 L=6e-07 W=6.81e-06 AD=2.9964e-12 AS=2.9964e-12 PD=1.45e-05 PS=1.45e-05 NRD=0.0646109 NRS=0.0646109 m=1 nf=1 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT nmos_1p2$$47119404 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
X0 1 2 3 4 nfet_05v0_I12 $T=-155 0 0 0 $X=-835 $Y=-620
.ENDS
***************************************
.SUBCKT ypass_gate vss 3 b d bb db ypass pcb vdd
** N=26 EP=9 IP=25 FDC=5
*.SEEDPROM
X2 bb b pcb vdd pfet_05v0_I09 $T=1240 50985 1 0 $X=200 $Y=43555
X3 bb db 3 vdd pfet_05v0_I09 $T=1250 43050 1 0 $X=210 $Y=35620
X4 b d 3 vdd pmos_1p2$$46889004 $T=1405 15300 1 0 $X=-25 $Y=7790
X5 b d ypass vss nmos_1p2$$47119404 $T=1405 24575 1 0 $X=260 $Y=17090
X6 bb db ypass vss nmos_1p2$$47119404 $T=1405 34595 1 0 $X=260 $Y=27110
.ENDS
***************************************
.SUBCKT mux821 1 2 3 4 5 6 7 8 9 13 14 15 16 17 18 19 20 21 22 23
+ 24 25 26 27 28 29 30 31 32 33 42 43 44 45 46 47 48
** N=86 EP=37 IP=165 FDC=48
*.SEEDPROM
M0 13 42 1 1 nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=1510 $Y=2370 $D=2
M1 16 43 1 1 nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=3750 $Y=2370 $D=2
M2 19 44 1 1 nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=7705 $Y=2370 $D=2
M3 22 45 1 1 nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=9945 $Y=2370 $D=2
M4 25 46 1 1 nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=13895 $Y=2370 $D=2
M5 28 47 1 1 nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=16135 $Y=2370 $D=2
M6 31 48 1 1 nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=20090 $Y=2370 $D=2
M7 2 9 1 1 nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=3.99e-13 PD=2.18e-06 PS=3.11e-06 NRD=0.912281 NRS=1.22807 m=1 nf=2 $X=22330 $Y=2370 $D=2
X10 5 3 7 8 pfet_05v0_I09 $T=23310 51440 1 0 $X=22270 $Y=44010
X11 5 6 2 8 pfet_05v0_I09 $T=23320 43505 1 0 $X=22280 $Y=36075
X12 3 4 2 8 pmos_1p2$$46889004 $T=23475 15755 1 0 $X=22045 $Y=8245
X13 3 4 9 1 nmos_1p2$$47119404 $T=23475 25030 1 0 $X=22330 $Y=17545
X14 5 6 9 1 nmos_1p2$$47119404 $T=23475 35050 1 0 $X=22330 $Y=27565
X15 1 13 15 4 14 6 42 7 8 ypass_gate $T=3490 455 1 180 $X=-1160 $Y=0
X16 1 16 18 4 17 6 43 7 8 ypass_gate $T=3490 455 0 0 $X=2385 $Y=0
X17 1 19 21 4 20 6 44 7 8 ypass_gate $T=9685 455 1 180 $X=5035 $Y=0
X18 1 22 24 4 23 6 45 7 8 ypass_gate $T=9685 455 0 0 $X=8580 $Y=0
X19 1 25 27 4 26 6 46 7 8 ypass_gate $T=15875 455 1 180 $X=11225 $Y=0
X20 1 28 30 4 29 6 47 7 8 ypass_gate $T=15875 455 0 0 $X=14770 $Y=0
X21 1 31 33 4 32 6 48 7 8 ypass_gate $T=22070 455 1 180 $X=17420 $Y=0
.ENDS
***************************************
.SUBCKT pfet_05v0_I12
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_05v0_I17
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_05v0_I10
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$202587180
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_05v0_I11
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pfet_05v0_I18 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pfet_05v0 L=6e-07 W=3.42e-06 AD=8.892e-13 AS=1.5048e-12 PD=4.46e-06 PS=8.6e-06 NRD=0.304094 NRS=0.51462 m=1 nf=2 $X=0 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT pfet_05v0_I13
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_1p2$$202595372
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$202586156
** N=3 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_1p2$$202596396
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pfet_05v0_I08
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_05v0_I13
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT wen_wm1 vss wep 3 4 5 6 7 8 9 10 11 12 13 men vdd wen GWEN 18 19
** N=43 EP=19 IP=113 FDC=31
M0 3 wen vss vss nfet_05v0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=1765 $Y=5060 $D=2
M1 6 men vss vss nfet_05v0 L=6e-07 W=1.37e-06 AD=3.562e-13 AS=6.028e-13 PD=1.89e-06 PS=3.62e-06 NRD=0.189781 NRS=0.321168 m=1 nf=1 $X=1765 $Y=8905 $D=2
M2 vss GWEN 3 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=2885 $Y=5060 $D=2
M3 vss vss 6 vss nfet_05v0 L=6e-07 W=1.37e-06 AD=6.028e-13 AS=3.562e-13 PD=3.62e-06 PS=1.89e-06 NRD=0.321168 NRS=0.189781 m=1 nf=1 $X=2885 $Y=8905 $D=2
M4 4 3 vss vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=5125 $Y=4650 $D=2
M5 5 6 vss vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=5125 $Y=9315 $D=2
M6 9 6 4 vss nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=7660 $Y=8385 $D=2
M7 7 10 vss vss nfet_05v0 L=6e-07 W=1.37e-06 AD=6.028e-13 AS=6.028e-13 PD=3.62e-06 PS=3.62e-06 NRD=0.321168 NRS=0.321168 m=1 nf=1 $X=8920 $Y=4240 $D=2
M8 11 5 9 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=9970 $Y=9700 $D=2
M9 vss 12 11 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=11090 $Y=9700 $D=2
M10 vss 9 12 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=13330 $Y=9700 $D=2
M11 13 12 vss vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=14450 $Y=9700 $D=2
M12 wep 7 vss vss nfet_05v0 L=6e-07 W=2.4e-06 AD=7.68e-13 AS=7.68e-13 PD=5.12e-06 PS=5.12e-06 NRD=1.2 NRS=1.2 m=1 nf=3 $X=12720 $Y=4810 $D=2
M13 vss 13 8 vss nfet_05v0 L=6e-07 W=1.37e-06 AD=6.028e-13 AS=6.028e-13 PD=3.62e-06 PS=3.62e-06 NRD=0.321168 NRS=0.321168 m=1 nf=1 $X=17810 $Y=9290 $D=2
M14 men 8 10 vss nfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.589e-12 PD=5.58e-06 PS=8.21e-06 NRD=0.229075 NRS=0.30837 m=1 nf=2 $X=20050 $Y=8385 $D=2
M15 vss 13 10 vss nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=22290 $Y=8385 $D=2
M16 18 wen vdd vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=1765 $Y=600 $D=8
M17 19 men vdd vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=1765 $Y=12055 $D=8
M18 3 GWEN 18 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=2885 $Y=600 $D=8
M19 6 vss 19 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=2885 $Y=12055 $D=8
M20 4 3 vdd vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=5125 $Y=600 $D=8
M21 5 6 vdd vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=5125 $Y=12055 $D=8
M22 9 5 4 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=1.17084e-12 AS=9.988e-13 PD=4.78598e-06 PS=5.42e-06 NRD=0.22722 NRS=0.193833 m=1 nf=1 $X=7660 $Y=12055 $D=8
M23 11 6 9 vdd pfet_05v0 L=6e-07 W=9.6e-07 AD=-6.87097e-13 AS=-6.48697e-13 PD=-2.78573e-06 PS=-2.70573e-06 NRD=-0.745548 NRS=-0.703882 m=1 nf=1 $X=9395 $Y=12055 $D=8
M24 vdd 12 11 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=1.14386e-12 PD=5.42e-06 PS=4.72975e-06 NRD=0.193833 NRS=0.221983 m=1 nf=1 $X=11090 $Y=12055 $D=8
M25 vdd 9 12 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=13330 $Y=12055 $D=8
M26 13 12 vdd vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=14450 $Y=12055 $D=8
M27 wep 7 vdd vdd pfet_05v0 L=6e-07 W=6e-06 AD=1.92e-12 AS=1.92e-12 PD=9.92e-06 PS=9.92e-06 NRD=0.48 NRS=0.48 m=1 nf=3 $X=12720 $Y=870 $D=8
M28 men 13 10 vdd pfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.58e-06 PS=1.084e-05 NRD=0.229075 NRS=0.387665 m=1 nf=2 $X=20050 $Y=12055 $D=8
X48 vdd 7 10 pfet_05v0_I18 $T=8920 2870 1 0 $X=7880 $Y=540
X49 vdd 8 13 pfet_05v0_I18 $T=16690 12625 0 0 $X=15650 $Y=12005
.ENDS
***************************************
.SUBCKT M1_PSUB$$44997676
** N=7 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pfet_05v0_I07
** N=6 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$46286892
** N=5 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_05v0_I06 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 nfet_05v0 L=6e-07 W=1.135e-05 AD=3.3596e-12 AS=3.3596e-12 PD=1.658e-05 PS=1.658e-05 NRD=0.651982 NRS=0.651982 m=1 nf=5 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT pfet_05v0_I16 1 2 3 4 5
** N=6 EP=5 IP=0 FDC=2
M0 2 4 1 2 pfet_05v0 L=6e-07 W=1.2e-06 AD=3.12e-13 AS=5.28e-13 PD=1.72e-06 PS=3.28e-06 NRD=0.216667 NRS=0.366667 m=1 nf=1 $X=0 $Y=0 $D=8
M1 3 5 2 2 pfet_05v0 L=6e-07 W=1.2e-06 AD=5.28e-13 AS=3.12e-13 PD=3.28e-06 PS=1.72e-06 NRD=0.366667 NRS=0.216667 m=1 nf=1 $X=1120 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nfet_05v0_I03 1 2 3 4 5
** N=5 EP=5 IP=0 FDC=2
M0 2 4 1 2 nfet_05v0 L=6e-07 W=6e-07 AD=1.56e-13 AS=2.64e-13 PD=1.12e-06 PS=2.08e-06 NRD=0.433333 NRS=0.733333 m=1 nf=1 $X=0 $Y=0 $D=2
M1 3 5 2 2 nfet_05v0 L=6e-07 W=6e-07 AD=2.64e-13 AS=1.56e-13 PD=2.08e-06 PS=1.12e-06 NRD=0.733333 NRS=0.433333 m=1 nf=1 $X=1120 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT pmos_1p2$$46285868
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$46281772
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pfet_05v0_I10
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_05v0_I05 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 nfet_05v0 L=6e-07 W=6e-07 AD=2.64e-13 AS=2.64e-13 PD=2.08e-06 PS=2.08e-06 NRD=0.733333 NRS=0.733333 m=1 nf=1 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT nfet_05v0_I21
** N=6 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sacntl_2 vss 2 pcb 4 5 6 7 8 9 10 11 18 19 20 21 22 23 24 25 26
+ se vdd men
** N=54 EP=23 IP=83 FDC=39
M0 2 11 vss vss nfet_05v0 L=6e-07 W=2.28e-06 AD=5.928e-13 AS=1.0032e-12 PD=3.32e-06 PS=6.32e-06 NRD=0.45614 NRS=0.77193 m=1 nf=2 $X=795 $Y=26115 $D=2
M1 4 men vss vss nfet_05v0 L=6e-07 W=5.7e-06 AD=1.6872e-12 AS=1.6872e-12 PD=9.8e-06 PS=9.8e-06 NRD=1.29825 NRS=1.29825 m=1 nf=5 $X=855 $Y=4275 $D=2
M2 vss 10 pcb vss nfet_05v0 L=6e-07 W=1.589e-05 AD=4.54e-12 AS=4.54e-12 PD=2.216e-05 PS=2.216e-05 NRD=0.881057 NRS=0.881057 m=1 nf=7 $X=1950 $Y=9235 $D=2
M3 5 4 vss vss nfet_05v0 L=6e-07 W=2.86e-06 AD=7.436e-13 AS=1.2584e-12 PD=3.38e-06 PS=6.6e-06 NRD=0.0909091 NRS=0.153846 m=1 nf=1 $X=10910 $Y=8645 $D=2
M4 6 11 5 vss nfet_05v0 L=6e-07 W=2.86e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=12030 $Y=8645 $D=2
M5 7 19 6 vss nfet_05v0 L=6e-07 W=2.86e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=13150 $Y=8645 $D=2
M6 8 19 7 vss nfet_05v0 L=6e-07 W=2.86e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=14270 $Y=8645 $D=2
M7 9 11 8 vss nfet_05v0 L=6e-07 W=2.86e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=15390 $Y=8645 $D=2
M8 vss 4 9 vss nfet_05v0 L=6e-07 W=2.86e-06 AD=1.2584e-12 AS=7.436e-13 PD=6.6e-06 PS=3.38e-06 NRD=0.153846 NRS=0.0909091 m=1 nf=1 $X=16510 $Y=8645 $D=2
M9 10 7 vss vss nfet_05v0 L=6e-07 W=5.22e-06 AD=1.3572e-12 AS=2.2968e-12 PD=6.26e-06 PS=1.22e-05 NRD=0.199234 NRS=0.337165 m=1 nf=2 $X=18750 $Y=8895 $D=2
M10 11 20 vss vss nfet_05v0 L=6e-07 W=1.44e-06 AD=6.336e-13 AS=6.336e-13 PD=3.76e-06 PS=3.76e-06 NRD=0.305556 NRS=0.305556 m=1 nf=1 $X=21255 $Y=4090 $D=2
M11 se 19 vss vss nfet_05v0 L=6e-07 W=9.08e-06 AD=2.3608e-12 AS=3.178e-12 PD=1.116e-05 PS=1.642e-05 NRD=0.45815 NRS=0.61674 m=1 nf=4 $X=19460 $Y=25030 $D=2
M12 2 11 vdd vdd pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=3.0008e-12 PD=7.86e-06 PS=1.54e-05 NRD=0.152493 NRS=0.258065 m=1 nf=2 $X=795 $Y=20945 $D=8
M13 4 men vdd vdd pfet_05v0 L=6e-07 W=1.135e-05 AD=3.3596e-12 AS=3.3596e-12 PD=1.658e-05 PS=1.658e-05 NRD=0.651982 NRS=0.651982 m=1 nf=5 $X=855 $Y=590 $D=8
M14 19 2 vdd vdd pfet_05v0 L=6e-07 W=6.81e-06 AD=1.7706e-12 AS=2.1792e-12 PD=8.37e-06 PS=1.1e-05 NRD=0.343612 NRS=0.422907 m=1 nf=3 $X=5370 $Y=20990 $D=8
M15 vdd 4 19 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=8730 $Y=20990 $D=8
M16 pcb 10 vdd vdd pfet_05v0 L=6e-07 W=4.09e-05 AD=1.0634e-11 AS=1.21023e-11 PD=4.61e-05 PS=4.6818e-05 NRD=0.635697 NRS=0.723472 m=1 nf=10 $X=830 $Y=14055 $D=8
M17 7 19 vdd vdd pfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.06e-06 PS=9.96e-06 NRD=0.0572687 NRS=0.0969163 m=1 nf=1 $X=14270 $Y=13710 $D=8
M18 vdd 11 7 vdd pfet_05v0 L=6e-07 W=4.54e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=15390 $Y=13710 $D=8
M19 7 4 vdd vdd pfet_05v0 L=6e-07 W=4.54e-06 AD=1.9976e-12 AS=1.1804e-12 PD=9.96e-06 PS=5.06e-06 NRD=0.0969163 NRS=0.0572687 m=1 nf=1 $X=16510 $Y=13710 $D=8
M20 vdd 25 26 vdd pfet_05v0 L=6e-07 W=1.2e-06 AD=5.28e-13 AS=5.28e-13 PD=3.28e-06 PS=3.28e-06 NRD=0.366667 NRS=0.366667 m=1 nf=1 $X=18950 $Y=1670 $D=8
M21 10 7 vdd vdd pfet_05v0 L=6e-07 W=1.362e-05 AD=4.3584e-12 AS=4.3584e-12 PD=2.008e-05 PS=2.008e-05 NRD=0.211454 NRS=0.211454 m=1 nf=3 $X=18750 $Y=13710 $D=8
M22 se 19 vdd vdd pfet_05v0 L=6e-07 W=2.72e-05 AD=7.072e-12 AS=8.0512e-12 PD=3.24e-05 PS=3.856e-05 NRD=0.955882 NRS=1.08824 m=1 nf=10 $X=12740 $Y=20450 $D=8
X23 vdd 11 20 pfet_05v0_I18 $T=21255 985 0 0 $X=20215 $Y=365
X27 vss 18 2 vss nfet_05v0_I06 $T=5370 25030 0 0 $X=4690 $Y=24410
X28 19 18 4 vss nfet_05v0_I06 $T=12415 25030 0 0 $X=11735 $Y=24410
X29 20 vdd 21 4 vss pfet_05v0_I16 $T=8080 1480 0 0 $X=7040 $Y=860
X30 22 vdd 23 21 22 pfet_05v0_I16 $T=11705 1480 0 0 $X=10665 $Y=860
X31 24 vdd 25 23 24 pfet_05v0_I16 $T=15325 1480 0 0 $X=14285 $Y=860
X32 20 vss 21 4 vss nfet_05v0_I03 $T=8080 4420 0 0 $X=7400 $Y=3800
X33 22 vss 23 21 22 nfet_05v0_I03 $T=11705 4420 0 0 $X=11025 $Y=3800
X34 24 vss 25 23 24 nfet_05v0_I03 $T=15325 4420 0 0 $X=14645 $Y=3800
X39 26 vss 25 vss nfet_05v0_I05 $T=18950 4420 0 0 $X=18270 $Y=3800
.ENDS
***************************************
.SUBCKT nfet_05v0_I09
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pfet_05v0_I14
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pfet_05v0_I04
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_05v0_I01
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT outbuf_oe q vss 3 4 5 15 16 17 18 vdd GWE se qp qn 24
** N=66 EP=15 IP=48 FDC=18
M0 vss 5 q vss nfet_05v0 L=6e-07 W=1.272e-05 AD=3.3072e-12 AS=4.0704e-12 PD=1.584e-05 PS=2.08e-05 NRD=0.735849 NRS=0.90566 m=1 nf=6 $X=395 $Y=2665 $D=2
M1 3 GWE vss vss nfet_05v0 L=6e-07 W=1.6e-06 AD=7.04e-13 AS=7.04e-13 PD=4.08e-06 PS=4.08e-06 NRD=0.275 NRS=0.275 m=1 nf=1 $X=8145 $Y=2720 $D=2
M2 17 3 vss vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=9.68e-13 PD=5.28e-06 PS=5.28e-06 NRD=0.2 NRS=0.2 m=1 nf=1 $X=10105 $Y=2700 $D=2
M3 vss 16 4 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=13175 $Y=12845 $D=2
M4 5 15 4 vss nfet_05v0 L=6e-07 W=6.81e-06 AD=2.1792e-12 AS=2.1792e-12 PD=1.1e-05 PS=1.1e-05 NRD=0.422907 NRS=0.422907 m=1 nf=3 $X=12455 $Y=2720 $D=2
M5 vss se 15 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=17045 $Y=4035 $D=2
M6 5 qn 18 vss nfet_05v0 L=6e-07 W=5.68e-06 AD=1.4768e-12 AS=1.988e-12 PD=6.72e-06 PS=9.92e-06 NRD=0.183099 NRS=0.246479 m=1 nf=2 $X=19905 $Y=1945 $D=2
M7 vss 3 18 vss nfet_05v0 L=6e-07 W=5.68e-06 AD=1.4768e-12 AS=1.988e-12 PD=6.72e-06 PS=9.92e-06 NRD=0.183099 NRS=0.246479 m=1 nf=2 $X=22145 $Y=1945 $D=2
M8 vdd 5 q vdd pfet_05v0 L=6e-07 W=2.268e-05 AD=5.8968e-12 AS=7.2576e-12 PD=2.58e-05 PS=3.408e-05 NRD=0.412698 NRS=0.507937 m=1 nf=6 $X=395 $Y=6190 $D=8
M9 3 GWE vdd vdd pfet_05v0 L=6e-07 W=4e-06 AD=1.76e-12 AS=1.76e-12 PD=8.88e-06 PS=8.88e-06 NRD=0.11 NRS=0.11 m=1 nf=1 $X=8145 $Y=6395 $D=8
M10 17 3 vdd vdd pfet_05v0 L=6e-07 W=4.5e-06 AD=1.98e-12 AS=1.98e-12 PD=9.88e-06 PS=9.88e-06 NRD=0.0977778 NRS=0.0977778 m=1 nf=1 $X=10105 $Y=6175 $D=8
M11 4 16 vdd vdd pfet_05v0 L=6e-07 W=2.28e-06 AD=5.928e-13 AS=1.24202e-12 PD=3.32e-06 PS=5.60564e-06 NRD=0.45614 NRS=0.955691 m=1 nf=2 $X=12055 $Y=10310 $D=8
M12 5 se 4 vdd pfet_05v0 L=6e-07 W=6.81e-06 AD=2.1792e-12 AS=2.1792e-12 PD=1.1e-05 PS=1.1e-05 NRD=0.422907 NRS=0.422907 m=1 nf=3 $X=12455 $Y=6395 $D=8
M13 16 5 vdd vdd pfet_05v0 L=6e-07 W=1.2e-06 AD=5.28e-13 AS=7.79385e-13 PD=3.28e-06 PS=2.57436e-06 NRD=0.366667 NRS=0.541239 m=1 nf=1 $X=15085 $Y=10250 $D=8
M14 vdd se 15 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=17045 $Y=7030 $D=8
M15 5 qp 24 vdd pfet_05v0 L=6e-07 W=1.134e-05 AD=2.9484e-12 AS=3.969e-12 PD=1.238e-05 PS=1.841e-05 NRD=0.0917108 NRS=0.123457 m=1 nf=2 $X=19680 $Y=6685 $D=8
M16 vdd 17 24 vdd pfet_05v0 L=6e-07 W=1.134e-05 AD=2.9484e-12 AS=3.969e-12 PD=1.238e-05 PS=1.841e-05 NRD=0.0917108 NRS=0.123457 m=1 nf=2 $X=21920 $Y=6685 $D=8
X22 vss 16 5 vss nfet_05v0_I05 $T=15150 13365 1 0 $X=14470 $Y=12145
.ENDS
***************************************
.SUBCKT pmos_1p2$$46887980 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pfet_05v0 L=6e-07 W=1.361e-05 AD=5.9884e-12 AS=5.9884e-12 PD=2.81e-05 PS=2.81e-05 NRD=0.0323292 NRS=0.0323292 m=1 nf=1 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT pmos_1p2$$46273580 1 2 3
** N=3 EP=3 IP=3 FDC=1
M0 2 3 1 1 pfet_05v0 L=6e-07 W=2.28e-06 AD=5.928e-13 AS=1.0032e-12 PD=3.32e-06 PS=6.32e-06 NRD=0.45614 NRS=0.77193 m=1 nf=2 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nmos_1p2$$46883884 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 nfet_05v0 L=6e-07 W=1.134e-05 AD=4.9896e-12 AS=4.9896e-12 PD=2.356e-05 PS=2.356e-05 NRD=0.0388007 NRS=0.0388007 m=1 nf=1 $X=-155 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT pfet_05v0_I03 1 2 3 4 5 6
** N=6 EP=6 IP=0 FDC=2
M0 2 4 1 6 pfet_05v0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=0 $Y=0 $D=8
M1 3 5 2 6 pfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=1120 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nfet_05v0_I02 1 2 3 4 5 6
** N=6 EP=6 IP=0 FDC=2
M0 2 4 1 6 nfet_05v0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=0 $Y=0 $D=2
M1 3 5 2 6 nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=1120 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT nmos_1p2$$46563372 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
M0 2 3 1 4 nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=-155 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT M1_NWELL_I01
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT din vss 2 3 4 d db 7 8 9 10 11 12 vdd datain men wep
** N=69 EP=16 IP=73 FDC=24
M0 2 4 vss vss nfet_05v0 L=6e-07 W=1.361e-05 AD=5.9884e-12 AS=5.9884e-12 PD=2.81e-05 PS=2.81e-05 NRD=0.0323292 NRS=0.0323292 m=1 nf=1 $X=260 $Y=10430 $D=2
M1 3 wep vss vss nfet_05v0 L=6e-07 W=1.14e-06 AD=7.866e-13 AS=7.923e-13 PD=3.66e-06 PS=3.67e-06 NRD=0.605263 NRS=0.609649 m=1 nf=1 $X=3600 $Y=38320 $D=2
M2 vss 10 4 vss nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=11165 $Y=8655 $D=2
M3 3 wep vdd vdd pfet_05v0 L=6e-07 W=2.97e-06 AD=1.13602e-12 AS=1.7523e-12 PD=4.5e-06 PS=8.3e-06 NRD=0.515152 NRS=0.794613 m=1 nf=2 $X=3025 $Y=35440 $D=8
M4 vdd 2 7 vdd pfet_05v0 L=6e-07 W=1.134e-05 AD=4.9896e-12 AS=4.9896e-12 PD=2.356e-05 PS=2.356e-05 NRD=0.0388007 NRS=0.0388007 m=1 nf=1 $X=6980 $Y=26220 $D=8
X5 4 vdd 10 vdd pfet_05v0_I09 $T=11165 455 0 0 $X=10125 $Y=-165
X6 d 2 3 vdd pmos_1p2$$46889004 $T=2655 26220 0 0 $X=1225 $Y=25510
X7 db 7 3 vdd pmos_1p2$$46889004 $T=4895 26220 0 0 $X=3465 $Y=25510
X9 vdd 2 4 pmos_1p2$$46887980 $T=415 26220 0 0 $X=-1015 $Y=25510
X10 vdd 12 men pmos_1p2$$46273580 $T=2920 7175 1 0 $X=1490 $Y=5355
X11 vdd 11 4 pmos_1p2$$46273580 $T=7060 8140 1 0 $X=5630 $Y=6320
X12 d 2 wep vss nmos_1p2$$46883884 $T=2655 12695 0 0 $X=1510 $Y=12010
X13 db 7 wep vss nmos_1p2$$46883884 $T=4895 12695 0 0 $X=3750 $Y=12010
X14 7 vss 2 vss nmos_1p2$$46883884 $T=7135 12695 0 0 $X=5990 $Y=12010
X15 8 vdd 9 datain 8 vdd pfet_05v0_I03 $T=2765 3195 0 0 $X=1725 $Y=2575
X16 9 10 11 men 12 vdd pfet_05v0_I03 $T=6905 3605 0 0 $X=5865 $Y=2985
X17 8 vss 9 datain 8 vss nfet_05v0_I02 $T=2765 1790 1 0 $X=2085 $Y=210
X18 9 10 11 12 men vss nfet_05v0_I02 $T=6905 725 0 0 $X=6225 $Y=105
X19 vss 12 men vss nmos_1p2$$46563372 $T=3470 9035 0 0 $X=2325 $Y=8350
X20 vss 11 4 vss nmos_1p2$$46563372 $T=7060 10495 1 0 $X=5915 $Y=8860
.ENDS
***************************************
.SUBCKT nmos_1p2$$46553132
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$46897196 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
M0 2 3 1 4 pfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.58e-06 PS=1.084e-05 NRD=0.229075 NRS=0.387665 m=1 nf=2 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT pmos_1p2$$46898220
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_1p2$$46551084
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sa 1 vss 3 4 qn qp 7 pcb vdd d db se
** N=105 EP=12 IP=47 FDC=27
M0 1 vss vss vss nfet_05v0 L=6e-07 W=3.41e-06 AD=8.866e-13 AS=1.5004e-12 PD=3.93e-06 PS=7.7e-06 NRD=0.0762463 NRS=0.129032 m=1 nf=1 $X=11660 $Y=16585 $D=2
M1 3 4 1 vss nfet_05v0 L=6e-07 W=3.41e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=12780 $Y=16585 $D=2
M2 4 1 3 vss nfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=1.7732e-12 PD=7.86e-06 PS=7.86e-06 NRD=0.152493 NRS=0.152493 m=1 nf=2 $X=13900 $Y=16585 $D=2
M3 7 4 vss vss nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=15170 $Y=8510 $D=2
M4 1 4 3 vss nfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=1.7732e-12 PD=7.86e-06 PS=7.86e-06 NRD=0.152493 NRS=0.152493 m=1 nf=2 $X=16140 $Y=16585 $D=2
M5 4 1 3 vss nfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=1.7732e-12 PD=7.86e-06 PS=7.86e-06 NRD=0.152493 NRS=0.152493 m=1 nf=2 $X=18380 $Y=16585 $D=2
M6 vss 7 qp vss nfet_05v0 L=6e-07 W=6.81e-06 AD=1.7706e-12 AS=2.1792e-12 PD=8.37e-06 PS=1.1e-05 NRD=0.343612 NRS=0.422907 m=1 nf=3 $X=17410 $Y=8510 $D=2
M7 1 4 3 vss nfet_05v0 L=6e-07 W=3.41e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=20620 $Y=16585 $D=2
M8 qn 1 vss vss nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=20770 $Y=8510 $D=2
M9 3 se vss vss nfet_05v0 L=6e-07 W=2.272e-05 AD=5.9072e-12 AS=6.9296e-12 PD=2.688e-05 PS=3.328e-05 NRD=0.732394 NRS=0.859155 m=1 nf=8 $X=12945 $Y=12550 $D=2
M10 vss vss 1 vss nfet_05v0 L=6e-07 W=3.41e-06 AD=1.5004e-12 AS=8.866e-13 PD=7.7e-06 PS=3.93e-06 NRD=0.129032 NRS=0.0762463 m=1 nf=1 $X=21740 $Y=16585 $D=2
M11 4 vdd vdd vdd pfet_05v0 L=6e-07 W=9.1e-07 AD=2.366e-13 AS=4.004e-13 PD=1.43e-06 PS=2.7e-06 NRD=0.285714 NRS=0.483516 m=1 nf=1 $X=13985 $Y=24010 $D=8
M12 vdd 1 4 vdd pfet_05v0 L=6e-07 W=9.1e-07 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=15105 $Y=24010 $D=8
M13 d pcb vdd vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=15755 $Y=30660 $D=8
M14 7 4 vdd vdd pfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.589e-12 PD=5.58e-06 PS=8.21e-06 NRD=0.229075 NRS=0.30837 m=1 nf=2 $X=15170 $Y=4385 $D=8
M15 4 pcb 1 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=16875 $Y=26330 $D=8
M16 db pcb d vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=16875 $Y=30660 $D=8
M17 1 4 vdd vdd pfet_05v0 L=6e-07 W=1.82e-06 AD=4.732e-13 AS=4.732e-13 PD=2.86e-06 PS=2.86e-06 NRD=0.571429 NRS=0.571429 m=1 nf=2 $X=16225 $Y=24010 $D=8
M18 vdd pcb db vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=17995 $Y=30660 $D=8
M19 4 1 vdd vdd pfet_05v0 L=6e-07 W=9.1e-07 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=18465 $Y=24010 $D=8
M20 qp 7 vdd vdd pfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.1804e-12 PD=5.58e-06 PS=5.58e-06 NRD=0.229075 NRS=0.229075 m=1 nf=2 $X=17410 $Y=4385 $D=8
M21 vdd vdd 4 vdd pfet_05v0 L=6e-07 W=9.1e-07 AD=4.004e-13 AS=2.366e-13 PD=2.7e-06 PS=1.43e-06 NRD=0.483516 NRS=0.285714 m=1 nf=1 $X=19585 $Y=24010 $D=8
M22 qn 1 vdd vdd pfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.589e-12 PD=5.58e-06 PS=8.21e-06 NRD=0.229075 NRS=0.30837 m=1 nf=2 $X=19650 $Y=4385 $D=8
X28 db 1 se vdd pmos_1p2$$46897196 $T=12475 26330 0 0 $X=11045 $Y=25620
X29 d 4 se vdd pmos_1p2$$46897196 $T=12475 30660 0 0 $X=11045 $Y=29950
X30 d 4 se vdd pmos_1p2$$46897196 $T=20400 26330 0 0 $X=18970 $Y=25620
X31 db 1 se vdd pmos_1p2$$46897196 $T=20400 30660 0 0 $X=18970 $Y=29950
.ENDS
***************************************
.SUBCKT saout_m2 1 VSS q datain pcb men VDD b[0] bb[0] WEN b[7] bb[7] bb[6] b[6] b[5] bb[5] bb[4] b[4] b[3] bb[3]
+ bb[2] b[2] b[1] bb[1] 54 GWE ypass[7] ypass[6] ypass[5] ypass[4] ypass[3] ypass[2] ypass[1] ypass[0] GWEN 78 79 80 81 82
+ 83 84
** N=135 EP=42 IP=161 FDC=187
*.SEEDPROM
X0 VSS 54 b[0] 74 bb[0] 77 pcb VDD ypass[0] 78 bb[7] b[7] 79 bb[6] b[6] 80 bb[5] b[5] 81 bb[4]
+ b[4] 82 bb[3] b[3] 83 bb[2] b[2] 84 bb[1] b[1] ypass[7] ypass[6] ypass[5] ypass[4] ypass[3] ypass[2] ypass[1]
+ mux821 $T=2765 83345 0 0 $X=-1345 $Y=83340
X1 VSS 1 86 89 90 87 92 96 91 97 93 94 95 men VDD WEN GWEN 85 88 wen_wm1 $T=1610 -16845 0 0 $X=100 $Y=-17385
X2 VSS 98 pcb 72 103 104 105 106 108 111 112 100 99 101 75 102 73 107 109 110
+ 76 VDD men
+ sacntl_2 $T=3160 150 0 0 $X=425 $Y=30
X3 q VSS 113 115 116 118 117 114 120 VDD GWE 76 134 135 119 outbuf_oe $T=3160 27580 0 0 $X=500 $Y=25785
X4 VSS 121 124 129 74 77 126 122 125 127 128 123 VDD datain men 1 din $T=1615 39060 0 0 $X=500 $Y=38775
X5 130 VSS 132 131 135 134 133 pcb VDD 74 77 76 sa $T=3160 43075 0 0 $X=1375 $Y=42095
.ENDS
***************************************
.SUBCKT 018SRAM_cell1_dummy 1 2 3 4 5 7
** N=9 EP=6 IP=0 FDC=4
*.SEEDPROM
M0 1 7 2 3 nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=180 $Y=260 $D=2
M1 3 5 1 3 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=1710 $D=2
M2 5 1 3 3 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=1710 $D=2
M3 5 7 4 3 nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=2220 $Y=260 $D=2
.ENDS
***************************************
.SUBCKT ICV_6 1 3 4 5 6 7 8 9 10 11
** N=15 EP=10 IP=18 FDC=8
*.SEEDPROM
X0 5 4 1 6 7 3 018SRAM_cell1_dummy $T=-3000 0 0 0 $X=-3340 $Y=-340
X1 9 8 1 10 11 3 018SRAM_cell1_dummy $T=0 0 0 0 $X=-340 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_13 1 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
** N=26 EP=17 IP=30 FDC=16
*.SEEDPROM
X0 1 1 3 4 5 6 7 8 9 10 ICV_6 $T=-6000 0 0 0 $X=-9340 $Y=-340
X1 1 1 11 12 13 14 15 16 17 18 ICV_6 $T=0 0 0 0 $X=-3340 $Y=-340
.ENDS
***************************************
.SUBCKT 018SRAM_strap1
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_14 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
** N=29 EP=17 IP=32 FDC=16
*.SEEDPROM
X0 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 ICV_13 $T=-3000 0 0 0 $X=-12340 $Y=-340
.ENDS
***************************************
.SUBCKT 018SRAM_cell1
** N=8 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT 018SRAM_cell1_2x 1 2 3 5 6 7 8 9 10
** N=12 EP=9 IP=16 FDC=8
*.SEEDPROM
M0 1 5 7 3 nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=180 $Y=3470 $D=2
M1 9 6 1 3 nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=180 $Y=4760 $D=2
M2 3 8 7 3 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=1840 $D=2
M3 3 10 9 3 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=6210 $D=2
M4 8 7 3 3 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=1840 $D=2
M5 10 9 3 3 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=6210 $D=2
M6 2 5 8 3 nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=2220 $Y=3470 $D=2
M7 10 6 2 3 nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=2220 $Y=4760 $D=2
.ENDS
***************************************
.SUBCKT ICV_31 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
** N=16 EP=15 IP=24 FDC=16
*.SEEDPROM
X0 5 6 2 3 4 9 11 10 12 018SRAM_cell1_2x $T=-3000 0 0 0 $X=-3340 $Y=-340
X1 7 8 2 3 4 13 15 14 16 018SRAM_cell1_2x $T=0 0 0 0 $X=-340 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_32 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
** N=26 EP=18 IP=32 FDC=40
*.SEEDPROM
M0 1 20 19 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=8060 $D=8
M1 1 24 23 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=9340 $D=8
M2 20 19 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=8060 $D=8
M3 24 23 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=9340 $D=8
M4 1 22 21 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=8060 $D=8
M5 1 26 25 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=9340 $D=8
M6 22 21 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=8060 $D=8
M7 26 25 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=9340 $D=8
X8 2 3 4 7 8 9 10 11 19 12 20 13 21 14 22 ICV_31 $T=0 0 0 0 $X=-3340 $Y=-340
X9 2 5 6 7 8 9 10 23 15 24 16 25 17 26 18 ICV_31 $T=0 9000 0 0 $X=-3340 $Y=8660
.ENDS
***************************************
.SUBCKT ICV_33 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
** N=30 EP=30 IP=36 FDC=80
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 15 16 17 18 19 20 21 22 ICV_32 $T=-6000 0 0 0 $X=-9340 $Y=-340
X1 1 2 3 4 5 6 11 12 13 14 23 24 25 26 27 28 29 30 ICV_32 $T=0 0 0 0 $X=-3340 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_34 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34
** N=50 EP=34 IP=60 FDC=176
*.SEEDPROM
M0 1 36 35 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-8370 $Y=17060 $D=8
M1 1 44 43 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-8370 $Y=18340 $D=8
M2 36 35 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-7230 $Y=17060 $D=8
M3 44 43 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-7230 $Y=18340 $D=8
M4 1 38 37 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-5370 $Y=17060 $D=8
M5 1 46 45 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-5370 $Y=18340 $D=8
M6 38 37 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-4230 $Y=17060 $D=8
M7 46 45 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-4230 $Y=18340 $D=8
M8 1 40 39 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=17060 $D=8
M9 1 48 47 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=18340 $D=8
M10 40 39 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=17060 $D=8
M11 48 47 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=18340 $D=8
M12 1 42 41 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=17060 $D=8
M13 1 50 49 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=18340 $D=8
M14 42 41 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=17060 $D=8
M15 50 49 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=18340 $D=8
X16 1 2 3 4 5 6 11 12 13 14 15 16 17 18 19 20 21 22 35 36
+ 37 38 23 24 25 26 39 40 41 42
+ ICV_33 $T=0 0 0 0 $X=-9340 $Y=-340
X17 1 2 7 8 9 10 11 12 13 14 15 16 17 18 43 44 45 46 27 28
+ 29 30 47 48 49 50 31 32 33 34
+ ICV_33 $T=0 18000 0 0 $X=-9340 $Y=17660
.ENDS
***************************************
.SUBCKT 018SRAM_strap1_2x
** N=10 EP=0 IP=12 FDC=0
.ENDS
***************************************
.SUBCKT ICV_10
** N=15 EP=0 IP=20 FDC=0
.ENDS
***************************************
.SUBCKT ICV_11
** N=19 EP=0 IP=24 FDC=0
.ENDS
***************************************
.SUBCKT ICV_27 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
** N=16 EP=15 IP=24 FDC=16
*.SEEDPROM
X0 5 6 2 3 4 9 11 10 12 018SRAM_cell1_2x $T=0 0 0 0 $X=-340 $Y=-340
X1 7 8 2 3 4 13 15 14 16 018SRAM_cell1_2x $T=3000 0 0 0 $X=2660 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_28 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
** N=26 EP=18 IP=32 FDC=40
*.SEEDPROM
M0 1 20 19 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=8060 $D=8
M1 1 24 23 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=9340 $D=8
M2 20 19 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=8060 $D=8
M3 24 23 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=9340 $D=8
M4 1 22 21 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=8060 $D=8
M5 1 26 25 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=9340 $D=8
M6 22 21 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=8060 $D=8
M7 26 25 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=9340 $D=8
X8 2 3 4 7 8 9 10 11 19 12 20 13 21 14 22 ICV_27 $T=0 0 0 0 $X=-340 $Y=-340
X9 2 5 6 7 8 9 10 23 15 24 16 25 17 26 18 ICV_27 $T=0 9000 0 0 $X=-340 $Y=8660
.ENDS
***************************************
.SUBCKT ICV_29 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
** N=30 EP=30 IP=36 FDC=80
*.SEEDPROM
X0 1 2 3 4 5 6 7 8 9 10 15 16 17 18 19 20 21 22 ICV_28 $T=0 0 0 0 $X=-340 $Y=-340
X1 1 2 3 4 5 6 11 12 13 14 23 24 25 26 27 28 29 30 ICV_28 $T=6000 0 0 0 $X=5660 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_30 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34
** N=50 EP=34 IP=60 FDC=176
*.SEEDPROM
M0 1 36 35 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=17060 $D=8
M1 1 44 43 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=18340 $D=8
M2 36 35 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=17060 $D=8
M3 44 43 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=18340 $D=8
M4 1 38 37 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=17060 $D=8
M5 1 46 45 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=18340 $D=8
M6 38 37 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=17060 $D=8
M7 46 45 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=18340 $D=8
M8 1 40 39 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=6630 $Y=17060 $D=8
M9 1 48 47 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=6630 $Y=18340 $D=8
M10 40 39 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=7770 $Y=17060 $D=8
M11 48 47 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=7770 $Y=18340 $D=8
M12 1 42 41 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=9630 $Y=17060 $D=8
M13 1 50 49 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=9630 $Y=18340 $D=8
M14 42 41 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=10770 $Y=17060 $D=8
M15 50 49 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=10770 $Y=18340 $D=8
X16 1 2 3 4 5 6 11 12 13 14 15 16 17 18 19 20 21 22 35 36
+ 37 38 23 24 25 26 39 40 41 42
+ ICV_29 $T=0 0 0 0 $X=-340 $Y=-340
X17 1 2 7 8 9 10 11 12 13 14 15 16 17 18 43 44 45 46 27 28
+ 29 30 47 48 49 50 31 32 33 34
+ ICV_29 $T=0 18000 0 0 $X=-340 $Y=17660
.ENDS
***************************************
.SUBCKT ICV_35 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32
+ 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52
+ 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72
+ 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92
+ 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112
+ 113 114 115 116 117 118
** N=118 EP=106 IP=168 FDC=704
*.SEEDPROM
X0 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 55 56
+ 57 58 59 60 61 62 63 64 65 66 67 68 69 70
+ ICV_34 $T=-42000 -4500 0 0 $X=-51340 $Y=-4840
X1 13 14 15 16 17 18 19 20 21 22 31 32 33 34 35 36 37 38 71 72
+ 73 74 75 76 77 78 79 80 81 82 83 84 85 86
+ ICV_34 $T=-30000 -4500 0 0 $X=-39340 $Y=-4840
X4 13 14 15 16 17 18 19 20 21 22 39 40 41 42 43 44 45 46 87 88
+ 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ ICV_30 $T=-12000 -4500 1 180 $X=-24340 $Y=-4840
X5 13 14 15 16 17 18 19 20 21 22 47 48 49 50 51 52 53 54 103 104
+ 105 106 107 108 109 110 111 112 113 114 115 116 117 118
+ ICV_30 $T=0 -4500 1 180 $X=-12340 $Y=-4840
.ENDS
***************************************
.SUBCKT ICV_15 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24
+ 25 26 27 28 29 30 31 32 33 34 35 36 37
** N=53 EP=33 IP=55 FDC=32
*.SEEDPROM
X0 4 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 ICV_13 $T=-15000 0 0 0 $X=-24340 $Y=-340
X1 4 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 ICV_14 $T=0 0 0 0 $X=-12340 $Y=-340
.ENDS
***************************************
.SUBCKT dcap_103_novia
** N=2 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_8
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_9
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT saout_R_m2 1 vss q pcb datain men vdd b[7] bb[7] WEN b[0] bb[0] bb[1] b[1] b[2] bb[2] bb[3] b[3] b[4] bb[4]
+ bb[5] b[5] b[6] bb[6] 54 GWE ypass[0] ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6] ypass[7] GWEN 74 75 76 77 78
+ 79 80
** N=131 EP=42 IP=161 FDC=187
*.SEEDPROM
X0 vss 54 b[7] 70 bb[7] 73 pcb vdd ypass[7] 74 bb[0] b[0] 75 bb[1] b[1] 76 bb[2] b[2] 77 bb[3]
+ b[3] 78 bb[4] b[4] 79 bb[5] b[5] 80 bb[6] b[6] ypass[0] ypass[1] ypass[2] ypass[3] ypass[4] ypass[5] ypass[6]
+ mux821 $T=2765 83310 0 0 $X=-1345 $Y=83305
X1 vss 1 82 85 86 83 88 92 87 93 89 90 91 men vdd WEN GWEN 81 84 wen_wm1 $T=1610 -16880 0 0 $X=100 $Y=-17420
X2 vss 94 pcb 68 99 100 101 102 104 107 108 96 95 97 71 98 69 103 105 106
+ 72 vdd men
+ sacntl_2 $T=3160 115 0 0 $X=425 $Y=-5
X3 q vss 109 111 112 114 113 110 116 vdd GWE 72 130 131 115 outbuf_oe $T=3160 27545 0 0 $X=500 $Y=25750
X4 vss 117 120 125 70 73 122 118 121 123 124 119 vdd datain men 1 din $T=1615 39025 0 0 $X=500 $Y=38740
X5 126 vss 128 127 131 130 129 pcb vdd 70 73 72 sa $T=3160 43040 0 0 $X=1375 $Y=42060
.ENDS
***************************************
.SUBCKT 018SRAM_strap1_bndry
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT 018SRAM_strap1_2x_bndry
** N=10 EP=0 IP=12 FDC=0
.ENDS
***************************************
.SUBCKT ICV_26
** N=15 EP=0 IP=20 FDC=0
.ENDS
***************************************
.SUBCKT 018SRAM_cell1_cutPC
** N=7 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_24 1 2 4 7 8 9 10
** N=10 EP=7 IP=14 FDC=8
*.SEEDPROM
M0 1 4 7 4 nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=180 $Y=-1030 $D=2
M1 9 4 1 4 nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=180 $Y=260 $D=2
M2 4 8 7 4 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=-2660 $D=2
M3 4 10 9 4 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=1710 $D=2
M4 8 7 4 4 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=-2660 $D=2
M5 10 9 4 4 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=1710 $D=2
M6 2 4 8 4 nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=2220 $Y=-1030 $D=2
M7 10 4 2 4 nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=2220 $Y=260 $D=2
.ENDS
***************************************
.SUBCKT ICV_25 1 2 7 8 9 10 11 12
** N=16 EP=8 IP=20 FDC=20
*.SEEDPROM
M0 1 14 13 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=-5440 $D=8
M1 1 16 15 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=-4160 $D=8
M2 14 13 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=-5440 $D=8
M3 16 15 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=-4160 $D=8
X4 7 8 2 9 10 13 14 ICV_24 $T=0 -9000 0 0 $X=-340 $Y=-13840
X5 7 8 2 15 16 11 12 ICV_24 $T=0 0 0 0 $X=-340 $Y=-4840
.ENDS
***************************************
.SUBCKT pmoscap_W2_5_477_R270
** N=26 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_19
** N=6 EP=0 IP=8 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_20
** N=10 EP=0 IP=12 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmoscap_W2_5_R270
** N=13 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT M1_PSUB_I05
** N=2827 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT M1_PSUB_I04
** N=2001 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pmos_1p2$$47513644
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_05v0_I19
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_1p2$$47641644
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pfet_05v0_I02
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT xpredec0_xa 2 3 13 29 30
** N=40 EP=5 IP=40 FDC=4
*.SEEDPROM
M0 40 29 2 3 nfet_05v0 L=6e-07 W=1.225e-05 AD=3.185e-12 AS=7.2275e-12 PD=1.277e-05 PS=2.568e-05 NRD=0.0212245 NRS=0.0481633 m=1 nf=1 $X=3255 $Y=2430 $D=2
M1 3 30 40 3 nfet_05v0 L=6e-07 W=1.225e-05 AD=7.28875e-12 AS=3.185e-12 PD=2.569e-05 PS=1.277e-05 NRD=0.0485714 NRS=0.0212245 m=1 nf=1 $X=4375 $Y=2430 $D=2
M2 2 29 13 13 pfet_05v0 L=6e-07 W=1.52e-05 AD=3.952e-12 AS=6.688e-12 PD=1.572e-05 PS=3.128e-05 NRD=0.0171053 NRS=0.0289474 m=1 nf=1 $X=3255 $Y=19540 $D=8
M3 13 30 2 13 pfet_05v0 L=6e-07 W=1.52e-05 AD=6.688e-12 AS=3.952e-12 PD=3.128e-05 PS=1.572e-05 NRD=0.0289474 NRS=0.0171053 m=1 nf=1 $X=4375 $Y=19540 $D=8
.ENDS
***************************************
.SUBCKT pmos_1p2$$47330348_161 1 2 3 4
** N=4 EP=4 IP=4 FDC=1
M0 2 3 1 4 pfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT alatch vss ab a vdd enb en
** N=16 EP=6 IP=24 FDC=8
M0 ab 12 vss vss nfet_05v0 L=6e-07 W=3.64e-06 AD=9.464e-13 AS=1.6016e-12 PD=4.68e-06 PS=9.04e-06 NRD=0.285714 NRS=0.483516 m=1 nf=2 $X=2590 $Y=1475 $D=2
M1 vss ab 11 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=3710 $Y=12935 $D=2
M2 a en 12 vss nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=6280 $Y=1020 $D=2
M3 11 enb 12 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=6280 $Y=12935 $D=2
M4 ab 12 vdd vdd pfet_05v0 L=6e-07 W=9.08e-06 AD=2.3608e-12 AS=3.9952e-12 PD=1.012e-05 PS=1.992e-05 NRD=0.114537 NRS=0.193833 m=1 nf=2 $X=2590 $Y=4695 $D=8
M5 a enb 12 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=6280 $Y=5895 $D=8
X10 11 vdd ab vdd pmos_1p2$$47330348_161 $T=3865 11540 1 0 $X=2435 $Y=9910
X11 12 11 en vdd pmos_1p2$$47330348_161 $T=6435 11540 1 0 $X=5005 $Y=9910
.ENDS
***************************************
.SUBCKT M1_PSUB$$47335468
** N=8 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT xpredec0_bot 1 2 3 8 9 10 11
** N=33 EP=7 IP=7 FDC=12
M0 2 33 1 1 nfet_05v0 L=6e-07 W=7.04e-06 AD=3.0976e-12 AS=3.0976e-12 PD=1.496e-05 PS=1.496e-05 NRD=0.0625 NRS=0.0625 m=1 nf=1 $X=3755 $Y=35615 $D=2
M1 3 2 1 1 nfet_05v0 L=6e-07 W=5.22e-06 AD=2.2968e-12 AS=2.2968e-12 PD=1.132e-05 PS=1.132e-05 NRD=0.0842912 NRS=0.0842912 m=1 nf=1 $X=6325 $Y=36010 $D=2
M2 2 33 8 8 pfet_05v0 L=6e-07 W=1.769e-05 AD=7.7836e-12 AS=7.7836e-12 PD=3.626e-05 PS=3.626e-05 NRD=0.0248728 NRS=0.0248728 m=1 nf=1 $X=3755 $Y=16320 $D=8
M3 3 2 8 8 pfet_05v0 L=6e-07 W=1.316e-05 AD=5.7904e-12 AS=5.7904e-12 PD=2.72e-05 PS=2.72e-05 NRD=0.0334347 NRS=0.0334347 m=1 nf=1 $X=6325 $Y=20855 $D=8
X4 1 33 9 8 11 10 alatch $T=350 -3160 0 0 $X=-100 $Y=-3165
.ENDS
***************************************
.SUBCKT xpredec0 vss vdd men clk A[1] A[0] x[3] x[2] x[1] x[0]
** N=99 EP=10 IP=158 FDC=56
M0 x[3] 90 vss vss nfet_05v0 L=6e-07 W=1.816e-05 AD=4.7216e-12 AS=5.5388e-12 PD=2.024e-05 PS=2.514e-05 NRD=0.229075 NRS=0.268722 m=1 nf=4 $X=260 $Y=50820 $D=2
M1 x[2] 92 vss vss nfet_05v0 L=6e-07 W=1.816e-05 AD=4.7216e-12 AS=4.7216e-12 PD=2.024e-05 PS=2.024e-05 NRD=0.229075 NRS=0.229075 m=1 nf=4 $X=4740 $Y=50820 $D=2
M2 x[1] 94 vss vss nfet_05v0 L=6e-07 W=1.816e-05 AD=4.7216e-12 AS=4.7216e-12 PD=2.024e-05 PS=2.024e-05 NRD=0.229075 NRS=0.229075 m=1 nf=4 $X=9220 $Y=50820 $D=2
M3 x[0] 96 vss vss nfet_05v0 L=6e-07 W=1.816e-05 AD=4.7216e-12 AS=5.5388e-12 PD=2.024e-05 PS=2.514e-05 NRD=0.229075 NRS=0.268722 m=1 nf=4 $X=13700 $Y=50820 $D=2
M4 17 men vss vss nfet_05v0 L=6e-07 W=1.37e-06 AD=3.562e-13 AS=6.028e-13 PD=1.89e-06 PS=3.62e-06 NRD=0.189781 NRS=0.321168 m=1 nf=1 $X=21630 $Y=51200 $D=2
M5 vss clk 17 vss nfet_05v0 L=6e-07 W=1.37e-06 AD=6.028e-13 AS=3.562e-13 PD=3.62e-06 PS=1.89e-06 NRD=0.321168 NRS=0.189781 m=1 nf=1 $X=22750 $Y=51200 $D=2
M6 x[3] 90 vdd vdd pfet_05v0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.38348e-11 PD=4.744e-05 PS=5.914e-05 NRD=0.0917108 NRS=0.107584 m=1 nf=4 $X=260 $Y=38080 $D=8
M7 x[2] 92 vdd vdd pfet_05v0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.744e-05 PS=4.744e-05 NRD=0.0917108 NRS=0.0917108 m=1 nf=4 $X=4740 $Y=38080 $D=8
M8 x[1] 94 vdd vdd pfet_05v0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.744e-05 PS=4.744e-05 NRD=0.0917108 NRS=0.0917108 m=1 nf=4 $X=9220 $Y=38080 $D=8
M9 x[0] 96 vdd vdd pfet_05v0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.38348e-11 PD=4.744e-05 PS=5.914e-05 NRD=0.0917108 NRS=0.107584 m=1 nf=4 $X=13700 $Y=38080 $D=8
M10 98 men vdd vdd pfet_05v0 L=6e-07 W=1.705e-06 AD=4.39037e-13 AS=1.01447e-12 PD=2.22e-06 PS=4.6e-06 NRD=0.151026 NRS=0.348974 m=1 nf=1 $X=21630 $Y=47525 $D=8
M11 17 clk 98 vdd pfet_05v0 L=6e-07 W=1.705e-06 AD=8.525e-15 AS=-8.525e-15 PD=1e-08 PS=-1e-08 NRD=0.00293255 NRS=-0.00293255 m=1 nf=1 $X=22745 $Y=47525 $D=8
M12 99 clk 17 vdd pfet_05v0 L=6e-07 W=1.705e-06 AD=-8.525e-15 AS=8.525e-15 PD=-1e-08 PS=1e-08 NRD=-0.00293255 NRS=0.00293255 m=1 nf=1 $X=23870 $Y=47525 $D=8
M13 vdd men 99 vdd pfet_05v0 L=6e-07 W=1.705e-06 AD=1.01447e-12 AS=4.39037e-13 PD=4.6e-06 PS=2.22e-06 NRD=0.348974 NRS=0.151026 m=1 nf=1 $X=24985 $Y=47525 $D=8
M14 18 17 vdd vdd pfet_05v0 L=6e-07 W=2.28e-06 AD=5.928e-13 AS=1.0032e-12 PD=3.32e-06 PS=6.32e-06 NRD=0.45614 NRS=0.77193 m=1 nf=2 $X=29010 $Y=47595 $D=8
X17 18 vss 17 vss nmos_1p2$$46563372 $T=29755 51180 0 0 $X=28610 $Y=50495
X18 90 vss vdd 30 31 xpredec0_xa $T=-2205 170 0 0 $X=-1440 $Y=-5
X19 92 vss vdd 30 32 xpredec0_xa $T=11165 170 1 180 $X=3000 $Y=-5
X20 94 vss vdd 33 31 xpredec0_xa $T=6755 170 0 0 $X=7520 $Y=-5
X21 96 vss vdd 33 32 xpredec0_xa $T=20125 170 1 180 $X=11960 $Y=-5
X22 vss 30 33 vdd A[1] 17 18 xpredec0_bot $T=18665 3160 0 0 $X=18135 $Y=-5
X23 vss 31 32 vdd A[0] 17 18 xpredec0_bot $T=27120 3160 0 0 $X=26590 $Y=-5
.ENDS
***************************************
.SUBCKT M1_PACTIVE_I03
** N=38 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pfet_05v0_I11
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_05v0_I14
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ypredec1_ys
** N=8 EP=0 IP=36 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_21 1 2 4 5 7 8
** N=8 EP=6 IP=10 FDC=4
*.SEEDPROM
M0 1 7 4 1 nfet_05v0 L=6e-07 W=2.724e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=3510 $Y=1700 $D=2
M1 8 5 1 1 nfet_05v0 L=6e-07 W=9.08e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=6870 $Y=1700 $D=2
M2 2 7 4 2 pfet_05v0 L=6e-07 W=6e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=3510 $Y=14855 $D=8
M3 8 5 2 2 pfet_05v0 L=6e-07 W=2e-05 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=6870 $Y=14855 $D=8
.ENDS
***************************************
.SUBCKT ICV_22 1 2 4 5 6 7 8 9 11 13
** N=14 EP=10 IP=16 FDC=12
*.SEEDPROM
M0 1 14 6 1 nfet_05v0 L=6e-07 W=2.724e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=9110 $Y=1700 $D=2
M1 12 7 1 1 nfet_05v0 L=6e-07 W=9.08e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=12470 $Y=1700 $D=2
M2 2 14 6 2 pfet_05v0 L=6e-07 W=6e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=9110 $Y=14855 $D=8
M3 12 7 2 2 pfet_05v0 L=6e-07 W=2e-05 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=12470 $Y=14855 $D=8
X4 1 2 4 5 11 14 ICV_21 $T=0 0 0 0 $X=-5 $Y=-5
X5 1 2 8 9 12 13 ICV_21 $T=11200 0 0 0 $X=11195 $Y=-5
.ENDS
***************************************
.SUBCKT nmos_1p2$$47514668
** N=4 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ypredec1_bot 1 2 3 10 11 12 13
** N=34 EP=7 IP=20 FDC=12
M0 2 30 1 1 nfet_05v0 L=6e-07 W=4.54e-06 AD=1.9976e-12 AS=1.9976e-12 PD=9.96e-06 PS=9.96e-06 NRD=0.0969163 NRS=0.0969163 m=1 nf=1 $X=3755 $Y=33350 $D=2
M1 3 2 1 1 nfet_05v0 L=6e-07 W=4.54e-06 AD=1.9976e-12 AS=1.9976e-12 PD=9.96e-06 PS=9.96e-06 NRD=0.0969163 NRS=0.0969163 m=1 nf=1 $X=6325 $Y=33350 $D=2
X2 10 2 30 pmos_1p2$$46887980 $T=3910 18340 0 0 $X=2480 $Y=17630
X3 10 3 2 pmos_1p2$$46887980 $T=6480 18340 0 0 $X=5050 $Y=17630
X4 1 30 11 10 13 12 alatch $T=350 -3160 0 0 $X=-100 $Y=-3165
.ENDS
***************************************
.SUBCKT pmos_1p2$$47821868
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$47820844
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ypredec1_xa
** N=29 EP=0 IP=36 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_23 1 2 5 8 9 10 11 12
** N=22 EP=8 IP=36 FDC=16
M0 20 10 13 1 nfet_05v0 L=6e-07 W=6.81e-06 AD=1.73655e-12 AS=4.05195e-12 PD=7.32e-06 PS=1.481e-05 NRD=0.0374449 NRS=0.0873715 m=1 nf=1 $X=-2370 $Y=-33035 $D=2
M1 19 9 20 1 nfet_05v0 L=6e-07 W=6.81e-06 AD=3.405e-14 AS=-3.405e-14 PD=1e-08 PS=-1e-08 NRD=0.000734214 NRS=-0.000734214 m=1 nf=1 $X=-1260 $Y=-33035 $D=2
M2 1 2 19 1 nfet_05v0 L=6e-07 W=6.81e-06 AD=3.405e-14 AS=-3.405e-14 PD=1e-08 PS=-1e-08 NRD=0.000734214 NRS=-0.000734214 m=1 nf=1 $X=-140 $Y=-33035 $D=2
M3 1 13 11 1 nfet_05v0 L=6e-07 W=6.81e-06 AD=1.7706e-12 AS=2.1792e-12 PD=8.37e-06 PS=1.1e-05 NRD=0.343612 NRS=0.422907 m=1 nf=3 $X=-2375 $Y=-2950 $D=2
M4 21 5 1 1 nfet_05v0 L=6e-07 W=6.81e-06 AD=-3.405e-14 AS=3.405e-14 PD=-1e-08 PS=1e-08 NRD=-0.000734214 NRS=0.000734214 m=1 nf=1 $X=990 $Y=-33035 $D=2
M5 22 9 21 1 nfet_05v0 L=6e-07 W=6.81e-06 AD=-3.405e-14 AS=3.405e-14 PD=-1e-08 PS=1e-08 NRD=-0.000734214 NRS=0.000734214 m=1 nf=1 $X=2110 $Y=-33035 $D=2
M6 16 10 22 1 nfet_05v0 L=6e-07 W=6.81e-06 AD=4.05195e-12 AS=1.73655e-12 PD=1.481e-05 PS=7.32e-06 NRD=0.0873715 NRS=0.0374449 m=1 nf=1 $X=3220 $Y=-33035 $D=2
M7 12 16 1 1 nfet_05v0 L=6e-07 W=6.81e-06 AD=2.1792e-12 AS=1.7706e-12 PD=1.1e-05 PS=8.37e-06 NRD=0.422907 NRS=0.343612 m=1 nf=3 $X=985 $Y=-2950 $D=2
M8 8 10 13 8 pfet_05v0 L=6e-07 W=5.67e-06 AD=1.4742e-12 AS=2.4948e-12 PD=6.19e-06 PS=1.222e-05 NRD=0.0458554 NRS=0.0776014 m=1 nf=1 $X=-2375 $Y=-19360 $D=8
M9 13 9 8 8 pfet_05v0 L=6e-07 W=5.67e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=-1255 $Y=-19360 $D=8
M10 8 2 13 8 pfet_05v0 L=6e-07 W=5.67e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=-135 $Y=-19360 $D=8
M11 8 13 11 8 pfet_05v0 L=6e-07 W=1.731e-05 AD=4.5006e-12 AS=5.5392e-12 PD=1.887e-05 PS=2.5e-05 NRD=0.135182 NRS=0.166378 m=1 nf=3 $X=-2375 $Y=-10125 $D=8
M12 16 5 8 8 pfet_05v0 L=6e-07 W=5.67e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=985 $Y=-19360 $D=8
M13 8 9 16 8 pfet_05v0 L=6e-07 W=5.67e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=2105 $Y=-19360 $D=8
M14 16 10 8 8 pfet_05v0 L=6e-07 W=5.67e-06 AD=2.4948e-12 AS=1.4742e-12 PD=1.222e-05 PS=6.19e-06 NRD=0.0776014 NRS=0.0458554 m=1 nf=1 $X=3225 $Y=-19360 $D=8
M15 12 16 8 8 pfet_05v0 L=6e-07 W=1.731e-05 AD=5.5392e-12 AS=4.5006e-12 PD=2.5e-05 PS=1.887e-05 NRD=0.166378 NRS=0.135182 m=1 nf=3 $X=985 $Y=-10125 $D=8
.ENDS
***************************************
.SUBCKT pmos_1p2$$47109164 1 2 3
** N=4 EP=3 IP=0 FDC=1
M0 2 3 1 1 pfet_05v0 L=6e-07 W=3.42e-06 AD=8.892e-13 AS=1.5048e-12 PD=4.46e-06 PS=8.6e-06 NRD=0.304094 NRS=0.51462 m=1 nf=2 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nmos_1p2$$47342636
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nfet_05v0_I07
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ypredec1 1 2 men clk ly[6] ly[7] ly[0] ly[1] ly[2] ly[3] ly[4] ly[5] ry[0] ry[1] ry[2] ry[3] ry[4] ry[5] ry[6] ry[7]
+ A[2] A[1] A[0]
** N=374 EP=23 IP=151 FDC=172
M0 367 358 1 1 nfet_05v0 L=6e-07 W=9.08e-06 AD=3.9952e-12 AS=3.9952e-12 PD=1.904e-05 PS=1.904e-05 NRD=0.0484581 NRS=0.0484581 m=1 nf=1 $X=2545 $Y=46970 $D=2
M1 1 371 ly[3] 1 nfet_05v0 L=6e-07 W=2.724e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=21585 $Y=46970 $D=2
M2 368 361 1 1 nfet_05v0 L=6e-07 W=9.08e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=24945 $Y=46970 $D=2
M3 188 189 1 1 nfet_05v0 L=6e-07 W=1.36e-06 AD=5.984e-13 AS=5.984e-13 PD=3.6e-06 PS=3.6e-06 NRD=0.323529 NRS=0.323529 m=1 nf=1 $X=31760 $Y=4985 $D=2
M4 189 clk 1 1 nfet_05v0 L=6e-07 W=1.91e-06 AD=4.966e-13 AS=8.404e-13 PD=2.43e-06 PS=4.7e-06 NRD=0.136126 NRS=0.230366 m=1 nf=1 $X=38610 $Y=5010 $D=2
M5 1 men 189 1 nfet_05v0 L=6e-07 W=1.91e-06 AD=8.404e-13 AS=4.966e-13 PD=4.7e-06 PS=2.43e-06 NRD=0.230366 NRS=0.136126 m=1 nf=1 $X=39730 $Y=5010 $D=2
M6 1 372 ly[7] 1 nfet_05v0 L=6e-07 W=2.724e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=43985 $Y=46970 $D=2
M7 369 358 1 1 nfet_05v0 L=6e-07 W=9.08e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=47345 $Y=46970 $D=2
M8 1 373 ry[3] 1 nfet_05v0 L=6e-07 W=2.724e-05 AD=7.0824e-12 AS=8.7168e-12 PD=2.88e-05 PS=3.824e-05 NRD=0.0859031 NRS=0.105727 m=1 nf=3 $X=66385 $Y=46970 $D=2
M9 370 361 1 1 nfet_05v0 L=6e-07 W=9.08e-06 AD=3.9952e-12 AS=2.3608e-12 PD=1.904e-05 PS=9.6e-06 NRD=0.0484581 NRS=0.0286344 m=1 nf=1 $X=69745 $Y=46970 $D=2
M10 1 374 ry[7] 1 nfet_05v0 L=6e-07 W=2.724e-05 AD=8.7168e-12 AS=8.7168e-12 PD=3.824e-05 PS=3.824e-05 NRD=0.105727 NRS=0.105727 m=1 nf=3 $X=88785 $Y=46970 $D=2
M11 367 358 2 2 pfet_05v0 L=6e-07 W=2e-05 AD=8.8e-12 AS=8.8e-12 PD=4.088e-05 PS=4.088e-05 NRD=0.022 NRS=0.022 m=1 nf=1 $X=2545 $Y=60125 $D=8
M12 2 371 ly[3] 2 pfet_05v0 L=6e-07 W=6e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=21585 $Y=60125 $D=8
M13 368 361 2 2 pfet_05v0 L=6e-07 W=2e-05 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=24945 $Y=60125 $D=8
M14 365 men 2 2 pfet_05v0 L=6e-07 W=2.275e-06 AD=5.915e-13 AS=1.35362e-12 PD=2.795e-06 PS=5.74e-06 NRD=0.114286 NRS=0.261538 m=1 nf=1 $X=36375 $Y=1335 $D=8
M15 189 clk 365 2 pfet_05v0 L=6e-07 W=2.275e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=37495 $Y=1335 $D=8
M16 366 clk 189 2 pfet_05v0 L=6e-07 W=2.275e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=38615 $Y=1335 $D=8
M17 2 men 366 2 pfet_05v0 L=6e-07 W=2.275e-06 AD=1.34225e-12 AS=5.915e-13 PD=5.73e-06 PS=2.795e-06 NRD=0.259341 NRS=0.114286 m=1 nf=1 $X=39735 $Y=1335 $D=8
M18 2 372 ly[7] 2 pfet_05v0 L=6e-07 W=6e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=43985 $Y=60125 $D=8
M19 369 358 2 2 pfet_05v0 L=6e-07 W=2e-05 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=47345 $Y=60125 $D=8
M20 2 373 ry[3] 2 pfet_05v0 L=6e-07 W=6e-05 AD=1.56e-11 AS=1.92e-11 PD=6.156e-05 PS=8.192e-05 NRD=0.039 NRS=0.048 m=1 nf=3 $X=66385 $Y=60125 $D=8
M21 370 361 2 2 pfet_05v0 L=6e-07 W=2e-05 AD=8.8e-12 AS=5.2e-12 PD=4.088e-05 PS=2.052e-05 NRD=0.022 NRS=0.013 m=1 nf=1 $X=69745 $Y=60125 $D=8
M22 2 374 ry[7] 2 pfet_05v0 L=6e-07 W=6e-05 AD=1.92e-11 AS=1.92e-11 PD=8.192e-05 PS=8.192e-05 NRD=0.048 NRS=0.048 m=1 nf=3 $X=88785 $Y=60125 $D=8
X23 1 2 ly[0] 357 ly[1] 359 ly[2] 360 367 371 ICV_22 $T=1275 45270 0 0 $X=1270 $Y=45265
X24 1 2 ly[4] 362 ly[5] 363 ly[6] 364 368 372 ICV_22 $T=23675 45270 0 0 $X=23670 $Y=45265
X25 1 2 ry[0] 357 ry[1] 359 ry[2] 360 369 373 ICV_22 $T=46075 45270 0 0 $X=46070 $Y=45265
X26 1 2 ry[4] 362 ry[5] 363 ry[6] 364 370 374 ICV_22 $T=68475 45270 0 0 $X=68470 $Y=45265
X27 1 190 191 2 A[2] 189 188 ypredec1_bot $T=1920 5135 0 0 $X=1820 $Y=1970
X28 1 192 193 2 A[1] 189 188 ypredec1_bot $T=10375 5135 0 0 $X=10275 $Y=1970
X29 1 194 195 2 A[0] 189 188 ypredec1_bot $T=18830 5135 0 0 $X=18730 $Y=1970
X30 1 195 194 2 192 190 363 364 ICV_23 $T=33645 42985 1 180 $X=28115 $Y=7365
X31 1 195 194 2 193 190 361 362 ICV_23 $T=41810 42985 1 180 $X=36280 $Y=7365
X32 1 195 194 2 192 191 359 360 ICV_23 $T=49980 42985 1 180 $X=44450 $Y=7365
X33 1 195 194 2 193 191 358 357 ICV_23 $T=58150 42985 1 180 $X=52620 $Y=7365
X34 2 188 189 pmos_1p2$$47109164 $T=32795 1405 1 180 $X=28795 $Y=720
.ENDS
***************************************
.SUBCKT pfet_05v0_I06
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT M1_POLY2_I01
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nfet_05v0_I15
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$49272876_R270 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pfet_05v0 L=6e-07 W=1.1e-05 AD=2.86e-12 AS=4.84e-12 PD=1.204e-05 PS=2.376e-05 NRD=0.0945455 NRS=0.16 m=1 nf=2 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT pfet_05v0_I17
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT xdec 1 2 men 6 vss 8 28 vdd
** N=103 EP=8 IP=41 FDC=6
*.SEEDPROM
M0 2 6 men vss nfet_05v0 L=6e-07 W=6.6e-06 AD=2.904e-12 AS=1.716e-12 PD=1.496e-05 PS=7.64e-06 NRD=0.266667 NRS=0.157576 m=1 nf=2 $X=37460 $Y=965 $D=2
M1 vss 8 6 vss nfet_05v0 L=6e-07 W=6.6e-07 AD=2.904e-13 AS=2.904e-13 PD=2.2e-06 PS=2.2e-06 NRD=0.666667 NRS=0.666667 m=1 nf=1 $X=45970 $Y=965 $D=2
M2 2 8 men vdd pfet_05v0 L=6e-07 W=6.6e-06 AD=2.904e-12 AS=1.716e-12 PD=1.496e-05 PS=7.64e-06 NRD=0.266667 NRS=0.157576 m=1 nf=2 $X=32185 $Y=965 $D=8
M3 vdd 8 6 vdd pfet_05v0 L=6e-07 W=1.59e-06 AD=6.996e-13 AS=6.996e-13 PD=4.06e-06 PS=4.06e-06 NRD=0.27673 NRS=0.27673 m=1 nf=1 $X=43020 $Y=965 $D=8
X12 vdd 1 2 pmos_1p2$$49272876_R270 $T=29780 1120 0 90 $X=23605 $Y=-360
X13 vdd 28 2 pmos_1p2$$49272876_R270 $T=91805 1120 1 90 $X=91120 $Y=-360
.ENDS
***************************************
.SUBCKT xdec8 vss xc xb xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] vdd 102 men 104 LWL[1] RWL[1] LWL[2] RWL[2] LWL[3] RWL[3] LWL[4]
+ RWL[4] LWL[5] RWL[5] LWL[6] RWL[6] 120 121 269 272 315 318
** N=334 EP=31 IP=608 FDC=126
*.SEEDPROM
M0 vss 274 273 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=16340 $Y=5740 $D=2
M1 vss 273 LWL[1] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=7020 $D=2
M2 vss 280 LWL[2] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=9260 $D=2
M3 280 281 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=16340 $Y=11660 $D=2
M4 vss 288 287 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=16340 $Y=14740 $D=2
M5 vss 287 LWL[3] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=16020 $D=2
M6 vss 294 LWL[4] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=18260 $D=2
M7 294 295 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=16340 $Y=20660 $D=2
M8 vss 302 301 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=16340 $Y=23740 $D=2
M9 vss 301 LWL[5] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=25020 $D=2
M10 vss 308 LWL[6] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=27260 $D=2
M11 308 309 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=16340 $Y=29660 $D=2
M12 vss 276 274 vss nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=46620 $Y=8140 $D=2
M13 281 283 vss vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=46620 $Y=9260 $D=2
M14 vss 290 288 vss nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=46620 $Y=17140 $D=2
M15 295 297 vss vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=46620 $Y=18260 $D=2
M16 vss 304 302 vss nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=46620 $Y=26140 $D=2
M17 309 311 vss vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=46620 $Y=27260 $D=2
M18 323 xa[1] 276 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=66460 $Y=5900 $D=2
M19 324 xb 323 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=66460 $Y=7020 $D=2
M20 vss xc 324 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=66460 $Y=8085 $D=2
M21 326 xc vss vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=66460 $Y=9315 $D=2
M22 325 xb 326 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=66460 $Y=10380 $D=2
M23 283 xa[2] 325 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=66460 $Y=11500 $D=2
M24 327 xa[3] 290 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=66460 $Y=14900 $D=2
M25 328 xb 327 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=66460 $Y=16020 $D=2
M26 vss xc 328 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=66460 $Y=17085 $D=2
M27 330 xc vss vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=66460 $Y=18315 $D=2
M28 329 xb 330 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=66460 $Y=19380 $D=2
M29 297 xa[4] 329 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=66460 $Y=20500 $D=2
M30 331 xa[5] 304 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=66460 $Y=23900 $D=2
M31 332 xb 331 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=66460 $Y=25020 $D=2
M32 vss xc 332 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=66460 $Y=26085 $D=2
M33 334 xc vss vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=66460 $Y=27315 $D=2
M34 333 xb 334 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=66460 $Y=28380 $D=2
M35 311 xa[6] 333 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=66460 $Y=29500 $D=2
M36 vss 274 279 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=100255 $Y=5740 $D=2
M37 vss 279 RWL[1] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=7020 $D=2
M38 vss 286 RWL[2] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=9260 $D=2
M39 286 281 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=100255 $Y=11660 $D=2
M40 vss 288 293 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=100255 $Y=14740 $D=2
M41 vss 293 RWL[3] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=16020 $D=2
M42 vss 300 RWL[4] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=18260 $D=2
M43 300 295 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=100255 $Y=20660 $D=2
M44 vss 302 307 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=100255 $Y=23740 $D=2
M45 vss 307 RWL[5] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=25020 $D=2
M46 vss 314 RWL[6] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=27260 $D=2
M47 314 309 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=100255 $Y=29660 $D=2
M48 LWL[1] 273 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=4665 $Y=5900 $D=8
M49 vdd 280 LWL[2] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=4665 $Y=9260 $D=8
M50 LWL[3] 287 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=4665 $Y=14900 $D=8
M51 vdd 294 LWL[4] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=4665 $Y=18260 $D=8
M52 LWL[5] 301 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=4665 $Y=23900 $D=8
M53 vdd 308 LWL[6] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=4665 $Y=27260 $D=8
M54 vdd xa[1] 276 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=71980 $Y=5900 $D=8
M55 276 xb vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=7020 $D=8
M56 vdd xc 276 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=8140 $D=8
M57 283 xc vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=9260 $D=8
M58 vdd xb 283 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=10380 $D=8
M59 283 xa[2] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=71980 $Y=11500 $D=8
M60 vdd xa[3] 290 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=71980 $Y=14900 $D=8
M61 290 xb vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=16020 $D=8
M62 vdd xc 290 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=17140 $D=8
M63 297 xc vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=18260 $D=8
M64 vdd xb 297 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=19380 $D=8
M65 297 xa[4] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=71980 $Y=20500 $D=8
M66 vdd xa[5] 304 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=71980 $Y=23900 $D=8
M67 304 xb vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=25020 $D=8
M68 vdd xc 304 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=26140 $D=8
M69 311 xc vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=27260 $D=8
M70 vdd xb 311 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=28380 $D=8
M71 311 xa[6] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=71980 $Y=29500 $D=8
M72 RWL[1] 279 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=106930 $Y=5900 $D=8
M73 vdd 286 RWL[2] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=106930 $Y=9260 $D=8
M74 RWL[3] 293 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=106930 $Y=14900 $D=8
M75 vdd 300 RWL[4] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=106930 $Y=18260 $D=8
M76 RWL[5] 307 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=106930 $Y=23900 $D=8
M77 vdd 314 RWL[6] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=106930 $Y=27260 $D=8
X78 269 102 men 270 vss 104 272 vdd xdec $T=5 4500 1 0 $X=0 $Y=-1140
X79 273 274 men 275 vss 276 279 vdd xdec $T=5 4500 0 0 $X=0 $Y=3385
X80 280 281 men 282 vss 283 286 vdd xdec $T=5 13500 1 0 $X=0 $Y=7860
X81 287 288 men 289 vss 290 293 vdd xdec $T=5 13500 0 0 $X=0 $Y=12385
X82 294 295 men 296 vss 297 300 vdd xdec $T=5 22500 1 0 $X=0 $Y=16860
X83 301 302 men 303 vss 304 307 vdd xdec $T=5 22500 0 0 $X=0 $Y=21385
X84 308 309 men 310 vss 311 314 vdd xdec $T=5 31500 1 0 $X=0 $Y=25860
X85 315 120 men 316 vss 121 318 vdd xdec $T=5 31500 0 0 $X=0 $Y=30385
.ENDS
***************************************
.SUBCKT xdec32 vss xc xb[3] xb[2] xb[1] xb[0] xa[7] xa[6] xa[5] xa[4] xa[3] xa[2] xa[1] xa[0] vdd LWL[0] LWL[1] LWL[2] LWL[3] LWL[4]
+ LWL[5] LWL[6] LWL[7] LWL[8] LWL[9] LWL[10] LWL[11] LWL[12] LWL[13] LWL[14] LWL[15] LWL[16] LWL[17] LWL[18] LWL[19] LWL[20] LWL[21] LWL[22] LWL[23] LWL[24]
+ LWL[25] LWL[26] LWL[27] LWL[28] LWL[29] LWL[30] LWL[31] RWL[1] RWL[2] RWL[3] RWL[4] RWL[5] RWL[6] RWL[7] RWL[8] RWL[9] RWL[10] RWL[11] RWL[12] RWL[13]
+ RWL[14] RWL[15] RWL[16] RWL[17] RWL[18] RWL[19] RWL[20] RWL[21] RWL[22] RWL[23] RWL[24] RWL[25] RWL[26] RWL[27] RWL[28] RWL[29] RWL[30] RWL[31] RWL[0] men
** N=357 EP=80 IP=544 FDC=608
M0 vss 326 LWL[0] vss nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=16340 $Y=260 $D=2
M1 326 310 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=16340 $Y=2660 $D=2
M2 vss 312 328 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=16340 $Y=32740 $D=2
M3 vss 328 LWL[7] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=34020 $D=2
M4 vss 330 LWL[8] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=36260 $D=2
M5 330 314 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=16340 $Y=38660 $D=2
M6 vss 316 332 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=16340 $Y=68740 $D=2
M7 vss 332 LWL[15] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=70020 $D=2
M8 vss 334 LWL[16] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=72260 $D=2
M9 334 318 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=16340 $Y=74660 $D=2
M10 vss 320 336 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=16340 $Y=104740 $D=2
M11 vss 336 LWL[23] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=106020 $D=2
M12 vss 338 LWL[24] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=16340 $Y=108260 $D=2
M13 338 322 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=16340 $Y=110660 $D=2
M14 vss 324 340 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=16340 $Y=140740 $D=2
M15 vss 340 LWL[31] vss nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=16340 $Y=142020 $D=2
M16 310 311 vss vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=9.68e-13 PD=5.28e-06 PS=5.28e-06 NRD=0.2 NRS=0.2 m=1 nf=1 $X=46620 $Y=260 $D=2
M17 vss 313 312 vss nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=46620 $Y=35140 $D=2
M18 314 315 vss vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=46620 $Y=36260 $D=2
M19 vss 317 316 vss nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=46620 $Y=71140 $D=2
M20 318 319 vss vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=46620 $Y=72260 $D=2
M21 vss 321 320 vss nfet_05v0 L=6e-07 W=2.2e-06 AD=5.72e-13 AS=9.68e-13 PD=2.72e-06 PS=5.28e-06 NRD=0.118182 NRS=0.2 m=1 nf=1 $X=46620 $Y=107140 $D=2
M22 322 323 vss vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=5.72e-13 PD=5.28e-06 PS=2.72e-06 NRD=0.2 NRS=0.118182 m=1 nf=1 $X=46620 $Y=108260 $D=2
M23 vss 325 324 vss nfet_05v0 L=6e-07 W=2.2e-06 AD=9.68e-13 AS=9.68e-13 PD=5.28e-06 PS=5.28e-06 NRD=0.2 NRS=0.2 m=1 nf=1 $X=46620 $Y=143140 $D=2
M24 343 xc vss vss nfet_05v0 L=6e-07 W=3.15e-06 AD=7.32375e-13 AS=2.079e-12 PD=3.615e-06 PS=7.62e-06 NRD=0.0738095 NRS=0.209524 m=1 nf=1 $X=66460 $Y=315 $D=2
M25 342 xb[0] 343 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=66460 $Y=1380 $D=2
M26 311 xa[0] 342 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=66460 $Y=2500 $D=2
M27 344 xa[7] 313 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=66460 $Y=32900 $D=2
M28 345 xb[0] 344 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=66460 $Y=34020 $D=2
M29 vss xc 345 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=66460 $Y=35085 $D=2
M30 347 xc vss vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=66460 $Y=36315 $D=2
M31 346 xb[1] 347 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=66460 $Y=37380 $D=2
M32 315 xa[0] 346 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=66460 $Y=38500 $D=2
M33 348 xa[7] 317 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=66460 $Y=68900 $D=2
M34 349 xb[1] 348 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=66460 $Y=70020 $D=2
M35 vss xc 349 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=66460 $Y=71085 $D=2
M36 351 xc vss vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=66460 $Y=72315 $D=2
M37 350 xb[2] 351 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=66460 $Y=73380 $D=2
M38 319 xa[0] 350 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=66460 $Y=74500 $D=2
M39 352 xa[7] 321 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=66460 $Y=104900 $D=2
M40 353 xb[2] 352 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=66460 $Y=106020 $D=2
M41 vss xc 353 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.59875e-13 AS=-2.59875e-13 PD=1.65e-07 PS=-1.65e-07 NRD=0.0261905 NRS=-0.0261905 m=1 nf=1 $X=66460 $Y=107085 $D=2
M42 355 xc vss vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-2.59875e-13 AS=2.59875e-13 PD=-1.65e-07 PS=1.65e-07 NRD=-0.0261905 NRS=0.0261905 m=1 nf=1 $X=66460 $Y=108315 $D=2
M43 354 xb[3] 355 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.6625e-14 AS=-8.6625e-14 PD=5.5e-08 PS=-5.5e-08 NRD=0.00873016 NRS=-0.00873016 m=1 nf=1 $X=66460 $Y=109380 $D=2
M44 323 xa[0] 354 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.25225e-12 AS=8.19e-13 PD=7.73e-06 PS=3.67e-06 NRD=0.226984 NRS=0.0825397 m=1 nf=1 $X=66460 $Y=110500 $D=2
M45 356 xa[7] 325 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=8.19e-13 AS=2.25225e-12 PD=3.67e-06 PS=7.73e-06 NRD=0.0825397 NRS=0.226984 m=1 nf=1 $X=66460 $Y=140900 $D=2
M46 357 xb[3] 356 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=-8.6625e-14 AS=8.6625e-14 PD=-5.5e-08 PS=5.5e-08 NRD=-0.00873016 NRS=0.00873016 m=1 nf=1 $X=66460 $Y=142020 $D=2
M47 vss xc 357 vss nfet_05v0 L=6e-07 W=3.15e-06 AD=2.079e-12 AS=7.32375e-13 PD=7.62e-06 PS=3.615e-06 NRD=0.209524 NRS=0.0738095 m=1 nf=1 $X=66460 $Y=143085 $D=2
M48 vss 327 RWL[0] vss nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=100255 $Y=260 $D=2
M49 327 310 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=100255 $Y=2660 $D=2
M50 vss 312 329 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=100255 $Y=32740 $D=2
M51 vss 329 RWL[7] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=34020 $D=2
M52 vss 331 RWL[8] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=36260 $D=2
M53 331 314 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=100255 $Y=38660 $D=2
M54 vss 316 333 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=100255 $Y=68740 $D=2
M55 vss 333 RWL[15] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=70020 $D=2
M56 vss 335 RWL[16] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=72260 $D=2
M57 335 318 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=100255 $Y=74660 $D=2
M58 vss 320 337 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=100255 $Y=104740 $D=2
M59 vss 337 RWL[23] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=106020 $D=2
M60 vss 339 RWL[24] vss nfet_05v0 L=6e-07 W=1e-05 AD=3e-12 AS=2.6e-12 PD=1.12e-05 PS=1.104e-05 NRD=0.12 NRS=0.104 m=1 nf=2 $X=100255 $Y=108260 $D=2
M61 339 322 vss vss nfet_05v0 L=6e-07 W=5e-06 AD=3.1e-12 AS=1.7e-12 PD=1.124e-05 PS=5.68e-06 NRD=0.124 NRS=0.068 m=1 nf=1 $X=100255 $Y=110660 $D=2
M62 vss 324 341 vss nfet_05v0 L=6e-07 W=5e-06 AD=1.7e-12 AS=3.1e-12 PD=5.68e-06 PS=1.124e-05 NRD=0.068 NRS=0.124 m=1 nf=1 $X=100255 $Y=140740 $D=2
M63 vss 341 RWL[31] vss nfet_05v0 L=6e-07 W=1e-05 AD=3.9e-12 AS=2.6e-12 PD=1.656e-05 PS=1.104e-05 NRD=0.156 NRS=0.104 m=1 nf=2 $X=100255 $Y=142020 $D=2
M64 vdd 326 LWL[0] vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=4665 $Y=260 $D=8
M65 LWL[7] 328 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=4665 $Y=32900 $D=8
M66 vdd 330 LWL[8] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=4665 $Y=36260 $D=8
M67 LWL[15] 332 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=4665 $Y=68900 $D=8
M68 vdd 334 LWL[16] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=4665 $Y=72260 $D=8
M69 LWL[23] 336 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=4665 $Y=104900 $D=8
M70 vdd 338 LWL[24] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=4665 $Y=108260 $D=8
M71 LWL[31] 340 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=4665 $Y=140900 $D=8
M72 311 xc vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=71980 $Y=260 $D=8
M73 vdd xb[0] 311 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=1380 $D=8
M74 311 xa[0] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=71980 $Y=2500 $D=8
M75 vdd xa[7] 313 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=71980 $Y=32900 $D=8
M76 313 xb[0] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=34020 $D=8
M77 vdd xc 313 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=35140 $D=8
M78 315 xc vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=36260 $D=8
M79 vdd xb[1] 315 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=37380 $D=8
M80 315 xa[0] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=71980 $Y=38500 $D=8
M81 vdd xa[7] 317 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=71980 $Y=68900 $D=8
M82 317 xb[1] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=70020 $D=8
M83 vdd xc 317 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=71140 $D=8
M84 319 xc vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=72260 $D=8
M85 vdd xb[2] 319 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=73380 $D=8
M86 319 xa[0] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=71980 $Y=74500 $D=8
M87 vdd xa[7] 321 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=71980 $Y=104900 $D=8
M88 321 xb[2] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=106020 $D=8
M89 vdd xc 321 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=107140 $D=8
M90 323 xc vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=108260 $D=8
M91 vdd xb[3] 323 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=109380 $D=8
M92 323 xa[0] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=71980 $Y=110500 $D=8
M93 vdd xa[7] 325 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=6.812e-13 AS=1.1528e-12 PD=3.14e-06 PS=6.12e-06 NRD=0.0992366 NRS=0.167939 m=1 nf=1 $X=71980 $Y=140900 $D=8
M94 325 xb[3] vdd vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=71980 $Y=142020 $D=8
M95 vdd xc 325 vdd pfet_05v0 L=6e-07 W=2.62e-06 AD=1.1528e-12 AS=6.812e-13 PD=6.12e-06 PS=3.14e-06 NRD=0.167939 NRS=0.0992366 m=1 nf=1 $X=71980 $Y=143140 $D=8
M96 vdd 327 RWL[0] vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=106930 $Y=260 $D=8
M97 RWL[7] 329 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=106930 $Y=32900 $D=8
M98 vdd 331 RWL[8] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=106930 $Y=36260 $D=8
M99 RWL[15] 333 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=106930 $Y=68900 $D=8
M100 vdd 335 RWL[16] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=106930 $Y=72260 $D=8
M101 RWL[23] 337 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=7.8e-12 PD=4.192e-05 PS=3.156e-05 NRD=0.096 NRS=0.078 m=1 nf=3 $X=106930 $Y=104900 $D=8
M102 vdd 339 RWL[24] vdd pfet_05v0 L=6e-07 W=3e-05 AD=7.8e-12 AS=9.6e-12 PD=3.156e-05 PS=4.192e-05 NRD=0.078 NRS=0.096 m=1 nf=3 $X=106930 $Y=108260 $D=8
M103 RWL[31] 341 vdd vdd pfet_05v0 L=6e-07 W=3e-05 AD=9.6e-12 AS=9.6e-12 PD=4.192e-05 PS=4.192e-05 NRD=0.096 NRS=0.096 m=1 nf=3 $X=106930 $Y=140900 $D=8
X104 vss xc xb[0] xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] vdd 310 men 311 LWL[1] RWL[1] LWL[2] RWL[2] LWL[3] RWL[3] LWL[4]
+ RWL[4] LWL[5] RWL[5] LWL[6] RWL[6] 312 313 326 327 328 329
+ xdec8 $T=0 0 0 0 $X=0 $Y=-1140
X105 vss xc xb[1] xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] vdd 314 men 315 LWL[9] RWL[9] LWL[10] RWL[10] LWL[11] RWL[11] LWL[12]
+ RWL[12] LWL[13] RWL[13] LWL[14] RWL[14] 316 317 330 331 332 333
+ xdec8 $T=0 36000 0 0 $X=0 $Y=34860
X106 vss xc xb[2] xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] vdd 318 men 319 LWL[17] RWL[17] LWL[18] RWL[18] LWL[19] RWL[19] LWL[20]
+ RWL[20] LWL[21] RWL[21] LWL[22] RWL[22] 320 321 334 335 336 337
+ xdec8 $T=0 72000 0 0 $X=0 $Y=70860
X107 vss xc xb[3] xa[1] xa[2] xa[3] xa[4] xa[5] xa[6] vdd 322 men 323 LWL[25] RWL[25] LWL[26] RWL[26] LWL[27] RWL[27] LWL[28]
+ RWL[28] LWL[29] RWL[29] LWL[30] RWL[30] 324 325 338 339 340 341
+ xdec8 $T=0 108000 0 0 $X=0 $Y=106860
.ENDS
***************************************
.SUBCKT M1_NWELL$$204218412
** N=49 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT nfet_05v0_I18 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 2 nfet_05v0 L=6e-07 W=1.011e-05 AD=4.4484e-12 AS=4.4484e-12 PD=2.11e-05 PS=2.11e-05 NRD=0.0435213 NRS=0.0435213 m=1 nf=1 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT M1_PACTIVE$$204148780
** N=13 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT pmos_1p2$$204216364 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pfet_05v0 L=6e-07 W=2.526e-05 AD=6.5676e-12 AS=1.11144e-11 PD=2.63e-05 PS=5.228e-05 NRD=0.0411718 NRS=0.0696754 m=1 nf=2 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT pfet_05v0_I01 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 2 3 1 4 pfet_05v0 L=6e-07 W=6.59e-06 AD=2.8996e-12 AS=2.8996e-12 PD=1.406e-05 PS=1.406e-05 NRD=0.0667678 NRS=0.0667678 m=1 nf=1 $X=0 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nfet_05v0_I04 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 2 nfet_05v0 L=6e-07 W=2.64e-06 AD=1.1616e-12 AS=1.1616e-12 PD=6.16e-06 PS=6.16e-06 NRD=0.166667 NRS=0.166667 m=1 nf=1 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT pfet_05v0_I05 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pfet_05v0 L=6e-07 W=4.72e-05 AD=1.2272e-11 AS=1.39712e-11 PD=5.24e-05 PS=6.256e-05 NRD=0.550847 NRS=0.627119 m=1 nf=10 $X=0 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nfet_05v0_I20 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nfet_05v0 L=6e-07 W=1.92e-05 AD=4.992e-12 AS=5.6832e-12 PD=2.44e-05 PS=2.896e-05 NRD=1.35417 NRS=1.54167 m=1 nf=10 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT M1_PACTIVE_I02
** N=7 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT wen_v2 vss vdd wen clk IGWEN GWE
** N=50 EP=6 IP=93 FDC=30
M0 vss wen 28 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=2545 $Y=1065 $D=2
M1 11 wen vss vss nfet_05v0 L=6e-07 W=6e-06 AD=1.92e-12 AS=1.92e-12 PD=9.92e-06 PS=9.92e-06 NRD=0.48 NRS=0.48 m=1 nf=3 $X=1260 $Y=16070 $D=2
M2 29 clk vss vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=3665 $Y=1065 $D=2
M3 30 29 vss vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=5905 $Y=1475 $D=2
M4 33 29 28 vss nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=8440 $Y=545 $D=2
M5 34 30 33 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=10750 $Y=1860 $D=2
M6 vss 35 34 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=11870 $Y=1860 $D=2
M7 vss 33 35 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=14110 $Y=1860 $D=2
M8 15 35 vss vss nfet_05v0 L=6e-07 W=2.4e-06 AD=6.24e-13 AS=1.056e-12 PD=3.44e-06 PS=6.56e-06 NRD=0.433333 NRS=0.733333 m=1 nf=2 $X=16465 $Y=1620 $D=2
M9 15 30 31 vss nfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.58e-06 PS=1.084e-05 NRD=0.229075 NRS=0.387665 m=1 nf=2 $X=19750 $Y=545 $D=2
M10 32 29 31 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=2.496e-13 AS=4.224e-13 PD=1.48e-06 PS=2.8e-06 NRD=0.270833 NRS=0.458333 m=1 nf=1 $X=23090 $Y=1240 $D=2
M11 vss 19 32 vss nfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=2.496e-13 PD=2.8e-06 PS=1.48e-06 NRD=0.458333 NRS=0.270833 m=1 nf=1 $X=24210 $Y=1240 $D=2
M12 19 31 vss vss nfet_05v0 L=6e-07 W=6.23e-06 AD=1.78e-12 AS=1.78e-12 PD=1.112e-05 PS=1.112e-05 NRD=2.24719 NRS=2.24719 m=1 nf=7 $X=26535 $Y=1905 $D=2
M13 vdd wen 28 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=5.902e-13 AS=9.988e-13 PD=2.79e-06 PS=5.42e-06 NRD=0.114537 NRS=0.193833 m=1 nf=1 $X=2545 $Y=4215 $D=8
M14 29 clk vdd vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=5.902e-13 PD=5.42e-06 PS=2.79e-06 NRD=0.193833 NRS=0.114537 m=1 nf=1 $X=3665 $Y=4215 $D=8
M15 30 29 vdd vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=5905 $Y=4215 $D=8
M16 11 wen vdd vdd pfet_05v0 L=6e-07 W=1.488e-05 AD=3.8688e-12 AS=4.7616e-12 PD=1.8e-05 PS=2.368e-05 NRD=0.629032 NRS=0.774194 m=1 nf=6 $X=1260 $Y=9420 $D=8
M17 33 30 28 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=1.17422e-12 AS=9.988e-13 PD=4.793e-06 PS=5.42e-06 NRD=0.227875 NRS=0.193833 m=1 nf=1 $X=8440 $Y=4215 $D=8
M18 34 29 33 vdd pfet_05v0 L=6e-07 W=9.6e-07 AD=-6.91897e-13 AS=-6.43897e-13 PD=-2.79573e-06 PS=-2.69573e-06 NRD=-0.750757 NRS=-0.698673 m=1 nf=1 $X=10180 $Y=4215 $D=8
M19 vdd 35 34 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=1.14048e-12 PD=5.42e-06 PS=4.72272e-06 NRD=0.193833 NRS=0.221328 m=1 nf=1 $X=11870 $Y=4215 $D=8
M20 vdd 33 35 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=14110 $Y=4215 $D=8
M21 15 35 vdd vdd pfet_05v0 L=6e-07 W=5.68e-06 AD=1.4768e-12 AS=2.4992e-12 PD=6.72e-06 PS=1.312e-05 NRD=0.183099 NRS=0.309859 m=1 nf=2 $X=16465 $Y=4215 $D=8
M22 15 29 31 vdd pfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=2.13253e-12 PD=5.58e-06 PS=1.01287e-05 NRD=0.229075 NRS=0.413851 m=1 nf=2 $X=19750 $Y=4215 $D=8
M23 32 30 31 vdd pfet_05v0 L=6e-07 W=9.6e-07 AD=-6.59976e-13 AS=-6.40776e-13 PD=-2.72923e-06 PS=-2.68923e-06 NRD=-0.71612 NRS=-0.695287 m=1 nf=1 $X=22550 $Y=5525 $D=8
M24 vdd 19 32 vdd pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=1.12024e-12 PD=5.42e-06 PS=4.68056e-06 NRD=0.193833 NRS=0.2174 m=1 nf=1 $X=24210 $Y=4215 $D=8
M25 19 31 vdd vdd pfet_05v0 L=6e-07 W=1.54e-05 AD=4.4e-12 AS=4.4e-12 PD=2.16e-05 PS=2.16e-05 NRD=0.909091 NRS=0.909091 m=1 nf=7 $X=26535 $Y=4215 $D=8
X46 vdd IGWEN 11 pfet_05v0_I05 $T=10115 9420 0 0 $X=9075 $Y=8800
X47 vdd GWE 19 pfet_05v0_I05 $T=23345 9420 0 0 $X=22305 $Y=8800
X48 vss IGWEN 11 nfet_05v0_I20 $T=10115 16070 0 0 $X=9435 $Y=15450
X49 vss GWE 19 nfet_05v0_I20 $T=23345 16070 0 0 $X=22665 $Y=15450
.ENDS
***************************************
.SUBCKT pmos_1p2$$47512620
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT xpredec1_xa
** N=29 EP=0 IP=36 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$47337516 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pfet_05v0 L=6e-07 W=1.633e-05 AD=7.1852e-12 AS=7.1852e-12 PD=3.354e-05 PS=3.354e-05 NRD=0.0269443 NRS=0.0269443 m=1 nf=1 $X=-155 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nmos_1p2$$47336492 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nfet_05v0 L=6e-07 W=6.58e-06 AD=2.8952e-12 AS=2.8952e-12 PD=1.404e-05 PS=1.404e-05 NRD=0.0668693 NRS=0.0668693 m=1 nf=1 $X=-155 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT xpredec1_bot 1 2 3 10 11 12 13
** N=32 EP=7 IP=19 FDC=12
X0 1 32 11 10 13 12 alatch $T=350 -3160 0 0 $X=-100 $Y=-3165
X2 10 2 32 pmos_1p2$$47337516 $T=3910 18340 0 0 $X=2480 $Y=17635
X3 10 3 2 pmos_1p2$$47337516 $T=6480 18340 0 0 $X=5050 $Y=17635
X4 1 2 32 nmos_1p2$$47336492 $T=3910 36070 0 0 $X=2765 $Y=35385
X5 1 3 2 nmos_1p2$$47336492 $T=6480 36070 0 0 $X=5335 $Y=35385
.ENDS
***************************************
.SUBCKT xpredec1 vss men vdd clk A[2] A[1] A[0] x[7] x[6] x[5] x[4] x[3] x[2] x[1] x[0]
** N=91 EP=15 IP=199 FDC=108
M0 77 18 51 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=3.2435e-12 AS=7.36025e-12 PD=1.2995e-05 PS=2.613e-05 NRD=0.0208417 NRS=0.0472946 m=1 nf=1 $X=1700 $Y=2310 $D=2
M1 76 19 77 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=2820 $Y=2310 $D=2
M2 vss 20 76 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=3940 $Y=2310 $D=2
M3 vss 51 x[7] vss nfet_05v0 L=6e-07 W=1.362e-05 AD=3.5412e-12 AS=4.3584e-12 PD=1.518e-05 PS=2.008e-05 NRD=0.171806 NRS=0.211454 m=1 nf=3 $X=1700 $Y=48000 $D=2
M4 78 21 vss vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=5060 $Y=2310 $D=2
M5 79 19 78 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=6180 $Y=2310 $D=2
M6 54 18 79 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=7.36025e-12 AS=3.2435e-12 PD=2.613e-05 PS=1.2995e-05 NRD=0.0472946 NRS=0.0208417 m=1 nf=1 $X=7300 $Y=2310 $D=2
M7 x[6] 54 vss vss nfet_05v0 L=6e-07 W=1.362e-05 AD=4.3584e-12 AS=3.5412e-12 PD=2.008e-05 PS=1.518e-05 NRD=0.211454 NRS=0.171806 m=1 nf=3 $X=5060 $Y=48000 $D=2
M8 81 18 57 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=3.2435e-12 AS=7.36025e-12 PD=1.2995e-05 PS=2.613e-05 NRD=0.0208417 NRS=0.0472946 m=1 nf=1 $X=9870 $Y=2310 $D=2
M9 80 22 81 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=10990 $Y=2310 $D=2
M10 vss 20 80 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=12110 $Y=2310 $D=2
M11 vss 57 x[5] vss nfet_05v0 L=6e-07 W=1.362e-05 AD=3.5412e-12 AS=4.3584e-12 PD=1.518e-05 PS=2.008e-05 NRD=0.171806 NRS=0.211454 m=1 nf=3 $X=9870 $Y=48000 $D=2
M12 82 21 vss vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=13230 $Y=2310 $D=2
M13 83 22 82 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=14350 $Y=2310 $D=2
M14 60 18 83 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=7.36025e-12 AS=3.2435e-12 PD=2.613e-05 PS=1.2995e-05 NRD=0.0472946 NRS=0.0208417 m=1 nf=1 $X=15470 $Y=2310 $D=2
M15 x[4] 60 vss vss nfet_05v0 L=6e-07 W=1.362e-05 AD=4.3584e-12 AS=3.5412e-12 PD=2.008e-05 PS=1.518e-05 NRD=0.211454 NRS=0.171806 m=1 nf=3 $X=13230 $Y=48000 $D=2
M16 85 23 63 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=3.2435e-12 AS=7.36025e-12 PD=1.2995e-05 PS=2.613e-05 NRD=0.0208417 NRS=0.0472946 m=1 nf=1 $X=18035 $Y=2310 $D=2
M17 84 19 85 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=19155 $Y=2310 $D=2
M18 vss 20 84 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=20275 $Y=2310 $D=2
M19 vss 63 x[3] vss nfet_05v0 L=6e-07 W=1.362e-05 AD=3.5412e-12 AS=4.3584e-12 PD=1.518e-05 PS=2.008e-05 NRD=0.171806 NRS=0.211454 m=1 nf=3 $X=18035 $Y=48000 $D=2
M20 86 21 vss vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=21395 $Y=2310 $D=2
M21 87 19 86 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=22515 $Y=2310 $D=2
M22 66 23 87 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=7.36025e-12 AS=3.2435e-12 PD=2.613e-05 PS=1.2995e-05 NRD=0.0472946 NRS=0.0208417 m=1 nf=1 $X=23635 $Y=2310 $D=2
M23 x[2] 66 vss vss nfet_05v0 L=6e-07 W=1.362e-05 AD=4.3584e-12 AS=3.5412e-12 PD=2.008e-05 PS=1.518e-05 NRD=0.211454 NRS=0.171806 m=1 nf=3 $X=21395 $Y=48000 $D=2
M24 89 23 69 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=3.2435e-12 AS=7.36025e-12 PD=1.2995e-05 PS=2.613e-05 NRD=0.0208417 NRS=0.0472946 m=1 nf=1 $X=26205 $Y=2310 $D=2
M25 88 22 89 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=27325 $Y=2310 $D=2
M26 vss 20 88 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=28445 $Y=2310 $D=2
M27 vss 69 x[1] vss nfet_05v0 L=6e-07 W=1.362e-05 AD=3.5412e-12 AS=4.3584e-12 PD=1.518e-05 PS=2.008e-05 NRD=0.171806 NRS=0.211454 m=1 nf=3 $X=26205 $Y=48000 $D=2
M28 90 21 vss vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=29565 $Y=2310 $D=2
M29 91 22 90 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=30685 $Y=2310 $D=2
M30 72 23 91 vss nfet_05v0 L=6e-07 W=1.2475e-05 AD=7.36025e-12 AS=3.2435e-12 PD=2.613e-05 PS=1.2995e-05 NRD=0.0472946 NRS=0.0208417 m=1 nf=1 $X=31805 $Y=2310 $D=2
M31 x[0] 72 vss vss nfet_05v0 L=6e-07 W=1.362e-05 AD=4.3584e-12 AS=3.5412e-12 PD=2.008e-05 PS=1.518e-05 NRD=0.211454 NRS=0.171806 m=1 nf=3 $X=29565 $Y=48000 $D=2
M32 17 men vss vss nfet_05v0 L=6e-07 W=1.91e-06 AD=4.966e-13 AS=8.404e-13 PD=2.43e-06 PS=4.7e-06 NRD=0.136126 NRS=0.230366 m=1 nf=1 $X=37165 $Y=51200 $D=2
M33 vss clk 17 vss nfet_05v0 L=6e-07 W=1.91e-06 AD=8.404e-13 AS=4.966e-13 PD=4.7e-06 PS=2.43e-06 NRD=0.230366 NRS=0.136126 m=1 nf=1 $X=38285 $Y=51200 $D=2
M34 vss 17 16 vss nfet_05v0 L=6e-07 W=1.36e-06 AD=5.984e-13 AS=5.984e-13 PD=3.6e-06 PS=3.6e-06 NRD=0.323529 NRS=0.323529 m=1 nf=1 $X=45140 $Y=51180 $D=2
M35 vdd 18 51 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=2.7118e-12 AS=4.5892e-12 PD=1.095e-05 PS=2.174e-05 NRD=0.0249281 NRS=0.042186 m=1 nf=1 $X=1700 $Y=21650 $D=8
M36 51 19 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=2820 $Y=21650 $D=8
M37 vdd 20 51 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=3940 $Y=21650 $D=8
M38 vdd 51 x[7] vdd pfet_05v0 L=6e-07 W=3.402e-05 AD=8.8452e-12 AS=1.08864e-11 PD=3.558e-05 PS=4.728e-05 NRD=0.0687831 NRS=0.0846561 m=1 nf=3 $X=1700 $Y=35260 $D=8
M39 54 21 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=5060 $Y=21650 $D=8
M40 vdd 19 54 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=6180 $Y=21650 $D=8
M41 54 18 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=4.5892e-12 AS=2.7118e-12 PD=2.174e-05 PS=1.095e-05 NRD=0.042186 NRS=0.0249281 m=1 nf=1 $X=7300 $Y=21650 $D=8
M42 x[6] 54 vdd vdd pfet_05v0 L=6e-07 W=3.402e-05 AD=1.08864e-11 AS=8.8452e-12 PD=4.728e-05 PS=3.558e-05 NRD=0.0846561 NRS=0.0687831 m=1 nf=3 $X=5060 $Y=35260 $D=8
M43 vdd 18 57 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=2.7118e-12 AS=4.5892e-12 PD=1.095e-05 PS=2.174e-05 NRD=0.0249281 NRS=0.042186 m=1 nf=1 $X=9870 $Y=21650 $D=8
M44 57 22 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=10990 $Y=21650 $D=8
M45 vdd 20 57 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=12110 $Y=21650 $D=8
M46 vdd 57 x[5] vdd pfet_05v0 L=6e-07 W=3.402e-05 AD=8.8452e-12 AS=1.08864e-11 PD=3.558e-05 PS=4.728e-05 NRD=0.0687831 NRS=0.0846561 m=1 nf=3 $X=9870 $Y=35260 $D=8
M47 60 21 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=13230 $Y=21650 $D=8
M48 vdd 22 60 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=14350 $Y=21650 $D=8
M49 60 18 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=4.5892e-12 AS=2.7118e-12 PD=2.174e-05 PS=1.095e-05 NRD=0.042186 NRS=0.0249281 m=1 nf=1 $X=15470 $Y=21650 $D=8
M50 x[4] 60 vdd vdd pfet_05v0 L=6e-07 W=3.402e-05 AD=1.08864e-11 AS=8.8452e-12 PD=4.728e-05 PS=3.558e-05 NRD=0.0846561 NRS=0.0687831 m=1 nf=3 $X=13230 $Y=35260 $D=8
M51 vdd 23 63 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=2.7118e-12 AS=4.5892e-12 PD=1.095e-05 PS=2.174e-05 NRD=0.0249281 NRS=0.042186 m=1 nf=1 $X=18035 $Y=21650 $D=8
M52 63 19 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=19155 $Y=21650 $D=8
M53 vdd 20 63 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=20275 $Y=21650 $D=8
M54 vdd 63 x[3] vdd pfet_05v0 L=6e-07 W=3.402e-05 AD=8.8452e-12 AS=1.08864e-11 PD=3.558e-05 PS=4.728e-05 NRD=0.0687831 NRS=0.0846561 m=1 nf=3 $X=18035 $Y=35260 $D=8
M55 66 21 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=21395 $Y=21650 $D=8
M56 vdd 19 66 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=22515 $Y=21650 $D=8
M57 66 23 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=4.5892e-12 AS=2.7118e-12 PD=2.174e-05 PS=1.095e-05 NRD=0.042186 NRS=0.0249281 m=1 nf=1 $X=23635 $Y=21650 $D=8
M58 x[2] 66 vdd vdd pfet_05v0 L=6e-07 W=3.402e-05 AD=1.08864e-11 AS=8.8452e-12 PD=4.728e-05 PS=3.558e-05 NRD=0.0846561 NRS=0.0687831 m=1 nf=3 $X=21395 $Y=35260 $D=8
M59 vdd 23 69 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=2.7118e-12 AS=4.5892e-12 PD=1.095e-05 PS=2.174e-05 NRD=0.0249281 NRS=0.042186 m=1 nf=1 $X=26205 $Y=21650 $D=8
M60 69 22 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=27325 $Y=21650 $D=8
M61 vdd 20 69 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=28445 $Y=21650 $D=8
M62 vdd 69 x[1] vdd pfet_05v0 L=6e-07 W=3.402e-05 AD=8.8452e-12 AS=1.08864e-11 PD=3.558e-05 PS=4.728e-05 NRD=0.0687831 NRS=0.0846561 m=1 nf=3 $X=26205 $Y=35260 $D=8
M63 72 21 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=29565 $Y=21650 $D=8
M64 vdd 22 72 vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=30685 $Y=21650 $D=8
M65 72 23 vdd vdd pfet_05v0 L=6e-07 W=1.043e-05 AD=4.5892e-12 AS=2.7118e-12 PD=2.174e-05 PS=1.095e-05 NRD=0.042186 NRS=0.0249281 m=1 nf=1 $X=31805 $Y=21650 $D=8
M66 x[0] 72 vdd vdd pfet_05v0 L=6e-07 W=3.402e-05 AD=1.08864e-11 AS=8.8452e-12 PD=4.728e-05 PS=3.558e-05 NRD=0.0846561 NRS=0.0687831 m=1 nf=3 $X=29565 $Y=35260 $D=8
M67 74 men vdd vdd pfet_05v0 L=6e-07 W=2.275e-06 AD=5.915e-13 AS=1.35362e-12 PD=2.795e-06 PS=5.74e-06 NRD=0.114286 NRS=0.261538 m=1 nf=1 $X=37165 $Y=47525 $D=8
M68 17 clk 74 vdd pfet_05v0 L=6e-07 W=2.275e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=38285 $Y=47525 $D=8
M69 75 clk 17 vdd pfet_05v0 L=6e-07 W=2.275e-06 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=39405 $Y=47525 $D=8
M70 vdd men 75 vdd pfet_05v0 L=6e-07 W=2.275e-06 AD=1.35362e-12 AS=5.915e-13 PD=5.74e-06 PS=2.795e-06 NRD=0.261538 NRS=0.114286 m=1 nf=1 $X=40525 $Y=47525 $D=8
X71 vdd 16 17 pmos_1p2$$47109164 $T=44700 47595 0 0 $X=42105 $Y=46910
X83 vss 18 23 vdd A[2] 17 16 xpredec1_bot $T=34205 3160 0 0 $X=33675 $Y=-5
X84 vss 19 22 vdd A[1] 17 16 xpredec1_bot $T=42655 3160 0 0 $X=42125 $Y=-5
X85 vss 20 21 vdd A[0] 17 16 xpredec1_bot $T=51110 3160 0 0 $X=50580 $Y=-5
.ENDS
***************************************
.SUBCKT pfet_05v0_I15 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pfet_05v0 L=1.2e-06 W=9e-07 AD=3.96e-13 AS=3.96e-13 PD=2.68e-06 PS=2.68e-06 NRD=0.488889 NRS=0.488889 m=1 nf=1 $X=0 $Y=0 $D=8
.ENDS
***************************************
.SUBCKT nfet_05v0_I16 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nfet_05v0 L=1.2e-06 W=6e-07 AD=2.64e-13 AS=2.64e-13 PD=2.08e-06 PS=2.08e-06 NRD=0.733333 NRS=0.733333 m=1 nf=1 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT pmos_1p2$$48624684
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_1p2$$47815724
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT strapx2b_bndry
** N=10 EP=0 IP=12 FDC=0
.ENDS
***************************************
.SUBCKT ICV_17 8 11 12 13 14 15 16
** N=16 EP=7 IP=22 FDC=8
*.SEEDPROM
X0 11 12 8 8 8 13 15 14 16 018SRAM_cell1_2x $T=0 0 0 0 $X=-340 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_18 7 8 13 14 18 19 20 21
** N=25 EP=8 IP=32 FDC=20
*.SEEDPROM
M0 7 23 22 7 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=8060 $D=8
M1 7 25 24 7 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=9340 $D=8
M2 23 22 7 7 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=8060 $D=8
M3 25 24 7 7 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=9340 $D=8
X4 8 13 14 18 22 19 23 ICV_17 $T=0 0 0 0 $X=-3340 $Y=-340
X5 8 13 14 24 20 25 21 ICV_17 $T=0 9000 0 0 $X=-3340 $Y=8660
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
** N=16 EP=16 IP=24 FDC=20
*.SEEDPROM
M0 1 12 9 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=8060 $D=8
M1 1 15 13 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=9340 $D=8
M2 12 9 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=8060 $D=8
M3 15 13 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=9340 $D=8
X4 8 10 2 3 4 7 11 9 12 018SRAM_cell1_2x $T=0 0 0 0 $X=-340 $Y=-340
X5 8 10 2 5 6 13 15 14 16 018SRAM_cell1_2x $T=0 9000 0 0 $X=-340 $Y=8660
.ENDS
***************************************
.SUBCKT ICV_5 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28
** N=28 EP=28 IP=32 FDC=44
*.SEEDPROM
M0 1 20 15 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=17060 $D=8
M1 1 25 21 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=18340 $D=8
M2 20 15 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=17060 $D=8
M3 25 21 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=18340 $D=8
X4 1 2 3 4 5 6 11 12 13 16 17 18 14 15 19 20 ICV_4 $T=0 0 0 0 $X=-340 $Y=-340
X5 1 2 7 8 9 10 21 12 22 16 25 26 23 24 27 28 ICV_4 $T=0 18000 0 0 $X=-340 $Y=17660
.ENDS
***************************************
.SUBCKT Cell_array32x1 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
** N=100 EP=100 IP=112 FDC=188
*.SEEDPROM
M0 1 52 43 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=35060 $D=8
M1 1 61 53 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=36340 $D=8
M2 1 68 60 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=71060 $D=8
M3 1 77 69 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=72340 $D=8
M4 1 84 76 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=107060 $D=8
M5 1 93 85 1 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=108340 $D=8
M6 52 43 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=35060 $D=8
M7 61 53 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=36340 $D=8
M8 68 60 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=71060 $D=8
M9 77 69 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=72340 $D=8
M10 84 76 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=107060 $D=8
M11 93 85 1 1 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=108340 $D=8
X12 1 2 3 4 5 6 7 8 9 10 35 36 37 38 39 44 45 46 47 48
+ 40 41 42 43 49 50 51 52
+ ICV_5 $T=0 0 0 0 $X=-340 $Y=-340
X13 1 2 11 12 13 14 15 16 17 18 53 36 54 55 56 44 61 62 63 64
+ 57 58 59 60 65 66 67 68
+ ICV_5 $T=0 36000 0 0 $X=-340 $Y=35660
X14 1 2 19 20 21 22 23 24 25 26 69 36 70 71 72 44 77 78 79 80
+ 73 74 75 76 81 82 83 84
+ ICV_5 $T=0 72000 0 0 $X=-340 $Y=71660
X15 1 2 27 28 29 30 31 32 33 34 85 36 86 87 88 44 93 94 95 96
+ 89 90 91 92 97 98 99 100
+ ICV_5 $T=0 108000 0 0 $X=-340 $Y=107660
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 48
+ 80 112 144
** N=175 EP=43 IP=215 FDC=392
*.SEEDPROM
M0 2 111 79 2 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=143060 $D=8
M1 2 45 47 2 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=144340 $D=8
M2 111 79 2 2 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=143060 $D=8
M3 45 47 2 2 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=144340 $D=8
M4 2 175 143 2 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=143060 $D=8
M5 2 41 43 2 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=3630 $Y=144340 $D=8
M6 175 143 2 2 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=143060 $D=8
M7 41 43 2 2 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=4770 $Y=144340 $D=8
X8 1 3 40 41 42 43 44 45 46 47 ICV_6 $T=3000 148500 0 180 $X=-340 $Y=143660
X9 2 1 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 48 36 49 50 51 52
+ 53 54 55 37 80 81 82 83 84 85 86 87 56 57 58 59 60 61 62 63
+ 88 89 90 91 92 93 94 95 64 65 66 67 68 69 70 71 96 97 98 99
+ 100 101 102 103 72 73 74 75 76 77 78 79 104 105 106 107 108 109 110 111
+ Cell_array32x1 $T=0 0 0 0 $X=-340 $Y=-340
X10 2 1 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 112 38 113 114 115 116
+ 117 118 119 39 144 145 146 147 148 149 150 151 120 121 122 123 124 125 126 127
+ 152 153 154 155 156 157 158 159 128 129 130 131 132 133 134 135 160 161 162 163
+ 164 165 166 167 136 137 138 139 140 141 142 143 168 169 170 171 172 173 174 175
+ Cell_array32x1 $T=3000 0 0 0 $X=2660 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_12
** N=27 EP=0 IP=32 FDC=0
.ENDS
***************************************
.SUBCKT ICV_7 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 48
+ 80 112 144
** N=175 EP=43 IP=215 FDC=392
*.SEEDPROM
M0 2 111 79 2 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=143060 $D=8
M1 2 43 41 2 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=-2370 $Y=144340 $D=8
M2 111 79 2 2 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=143060 $D=8
M3 43 41 2 2 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=-1230 $Y=144340 $D=8
M4 2 175 143 2 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=143060 $D=8
M5 2 47 45 2 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=144340 $D=8
M6 175 143 2 2 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=143060 $D=8
M7 47 45 2 2 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=144340 $D=8
X8 1 3 40 41 42 43 44 45 46 47 ICV_6 $T=0 148500 1 0 $X=-3340 $Y=143660
X9 2 1 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 48 36 49 50 51 52
+ 53 54 55 37 80 81 82 83 84 85 86 87 56 57 58 59 60 61 62 63
+ 88 89 90 91 92 93 94 95 64 65 66 67 68 69 70 71 96 97 98 99
+ 100 101 102 103 72 73 74 75 76 77 78 79 104 105 106 107 108 109 110 111
+ Cell_array32x1 $T=-3000 0 0 0 $X=-3340 $Y=-340
X10 2 1 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 112 38 113 114 115 116
+ 117 118 119 39 144 145 146 147 148 149 150 151 120 121 122 123 124 125 126 127
+ 152 153 154 155 156 157 158 159 128 129 130 131 132 133 134 135 160 161 162 163
+ 164 165 166 167 136 137 138 139 140 141 142 143 168 169 170 171 172 173 174 175
+ Cell_array32x1 $T=0 0 0 0 $X=-340 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_3
** N=15 EP=0 IP=20 FDC=0
.ENDS
***************************************
.SUBCKT 018SRAM_cell1_dummy_R
** N=8 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_1 3 4 7 8 9 10
** N=12 EP=6 IP=16 FDC=4
*.SEEDPROM
M0 4 4 7 4 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=3560 $D=8
M1 4 4 9 4 pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=630 $Y=4840 $D=8
M2 8 3 4 4 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=3560 $D=8
M3 10 3 4 4 pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=1770 $Y=4840 $D=8
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 10 12 14 15
** N=19 EP=8 IP=24 FDC=16
*.SEEDPROM
M0 1 3 16 3 nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=180 $Y=7970 $D=2
M1 18 3 1 3 nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=180 $Y=9260 $D=2
M2 3 4 16 3 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=6340 $D=2
M3 3 4 18 3 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=630 $Y=10710 $D=2
M4 17 3 3 3 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=6340 $D=2
M5 19 3 3 3 nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=1770 $Y=10710 $D=2
M6 2 3 17 3 nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=2220 $Y=7970 $D=2
M7 19 3 2 3 nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=2220 $Y=9260 $D=2
X8 3 4 10 12 16 17 ICV_1 $T=0 0 0 0 $X=-340 $Y=-340
X9 3 4 18 19 14 15 ICV_1 $T=0 9000 0 0 $X=-340 $Y=8660
.ENDS
***************************************
.SUBCKT gf180mcu_fd_ip_sram__sram256x8m8wm1 A[7] A[6] A[5] A[4] A[3] A[2] A[1]
+ A[0] CEN CLK D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] GWEN Q[7] Q[6] Q[5]
+ Q[4] Q[3] Q[2] Q[1] Q[0] VDD VSS WEN[7] WEN[6] WEN[5] WEN[4] WEN[3] WEN[2]
+ WEN[1] WEN[0]
** N=5478 EP=37 IP=4140 FDC=16461
M0 4301 VSS 712 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=120390 $Y=176390 $D=2
M1 712 VSS 4303 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=120390 $Y=328100 $D=2
M2 VSS 4300 4301 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=120840 $Y=177840 $D=2
M3 VSS 4302 4303 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=120840 $Y=326470 $D=2
M4 4300 4301 VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=121980 $Y=177840 $D=2
M5 4302 4303 VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=121980 $Y=326470 $D=2
M6 4300 VSS 711 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=122430 $Y=176390 $D=2
M7 711 VSS 4302 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=122430 $Y=328100 $D=2
M8 2 VDD 1 VSS nfet_05v0 L=6e-07 W=6.59e-06 AD=2.8996e-12 AS=2.8996e-12 PD=1.406e-05 PS=1.406e-05 NRD=0.0667678 NRS=0.0667678 m=1 nf=1 $X=204815 $Y=327000 $D=2
M9 VSS 1 802 VSS nfet_05v0 L=6e-07 W=1.36e-06 AD=3.536e-13 AS=5.984e-13 PD=1.88e-06 PS=3.6e-06 NRD=0.191176 NRS=0.323529 m=1 nf=1 $X=233770 $Y=54135 $D=2
M10 802 CLK VSS VSS nfet_05v0 L=6e-07 W=1.36e-06 AD=5.984e-13 AS=3.536e-13 PD=3.6e-06 PS=1.88e-06 NRD=0.323529 NRS=0.191176 m=1 nf=1 $X=234890 $Y=54135 $D=2
M11 616 619 VSS VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=1.1804e-12 AS=1.9976e-12 PD=5.58e-06 PS=1.084e-05 NRD=0.229075 NRS=0.387665 m=1 nf=2 $X=242235 $Y=54135 $D=2
M12 281 808 VSS VSS nfet_05v0 L=1e-06 W=6e-07 AD=2.64e-13 AS=2.64e-13 PD=2.08e-06 PS=2.08e-06 NRD=0.733333 NRS=0.733333 m=1 nf=1 $X=243265 $Y=46010 $D=2
M13 CEN 802 619 VSS nfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=245925 $Y=54135 $D=2
M14 250 468 VSS VSS nfet_05v0 L=6e-07 W=4.99e-05 AD=1.47704e-11 AS=1.47704e-11 PD=6.284e-05 PS=6.284e-05 NRD=0.148297 NRS=0.148297 m=1 nf=5 $X=241995 $Y=72320 $D=2
M15 317 281 VSS VSS nfet_05v0 L=6e-07 W=7.5e-07 AD=3.3e-13 AS=3.3e-13 PD=2.38e-06 PS=2.38e-06 NRD=0.586667 NRS=0.586667 m=1 nf=1 $X=246495 $Y=46075 $D=2
M16 354 317 VSS VSS nfet_05v0 L=6e-07 W=3.02e-06 AD=1.3288e-12 AS=1.3288e-12 PD=6.92e-06 PS=6.92e-06 NRD=0.145695 NRS=0.145695 m=1 nf=1 $X=249065 $Y=46070 $D=2
M17 4728 354 VSS VSS nfet_05v0 L=6e-07 W=2.268e-05 AD=5.8968e-12 AS=1.34946e-11 PD=2.32e-05 PS=4.655e-05 NRD=0.0114638 NRS=0.0262346 m=1 nf=1 $X=256125 $Y=28435 $D=2
M18 4729 CLK 4728 VSS nfet_05v0 L=6e-07 W=2.268e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=257245 $Y=28435 $D=2
M19 445 616 4729 VSS nfet_05v0 L=6e-07 W=2.268e-05 AD=1.33812e-11 AS=5.8968e-12 PD=4.654e-05 PS=2.32e-05 NRD=0.0260141 NRS=0.0114638 m=1 nf=1 $X=258365 $Y=28435 $D=2
M20 4730 495 VSS VSS nfet_05v0 L=6e-07 W=1.8145e-05 AD=4.7177e-12 AS=1.07963e-11 PD=1.8665e-05 PS=3.748e-05 NRD=0.014329 NRS=0.0327914 m=1 nf=1 $X=262120 $Y=29545 $D=2
M21 468 445 4730 VSS nfet_05v0 L=6e-07 W=1.8145e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=263240 $Y=29545 $D=2
M22 4731 445 468 VSS nfet_05v0 L=6e-07 W=1.8145e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=264360 $Y=29545 $D=2
M23 VSS 495 4731 VSS nfet_05v0 L=6e-07 W=1.8145e-05 AD=1.07055e-11 AS=4.7177e-12 PD=3.747e-05 PS=1.8665e-05 NRD=0.0325158 NRS=0.014329 m=1 nf=1 $X=265480 $Y=29545 $D=2
M24 4732 468 VSS VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=1.16905e-12 AS=2.7013e-12 PD=5.055e-06 PS=1.027e-05 NRD=0.0567181 NRS=0.131057 m=1 nf=1 $X=268545 $Y=43150 $D=2
M25 495 607 4732 VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=2.27e-14 AS=-2.27e-14 PD=1e-08 PS=-1e-08 NRD=0.00110132 NRS=-0.00110132 m=1 nf=1 $X=269660 $Y=43150 $D=2
M26 4733 607 495 VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=-2.27e-14 AS=2.27e-14 PD=-1e-08 PS=1e-08 NRD=-0.00110132 NRS=0.00110132 m=1 nf=1 $X=270785 $Y=43150 $D=2
M27 VSS 468 4733 VSS nfet_05v0 L=6e-07 W=4.54e-06 AD=2.7013e-12 AS=1.16905e-12 PD=1.027e-05 PS=5.055e-06 NRD=0.131057 NRS=0.0567181 m=1 nf=1 $X=271900 $Y=43150 $D=2
M28 1 250 VSS VSS nfet_05v0 L=6e-07 W=0.0001474 AD=3.8324e-11 AS=4.09772e-11 PD=0.0001578 PS=0.00017326 NRD=0.705563 NRS=0.75441 m=1 nf=20 $X=253180 $Y=76320 $D=2
M29 4305 VSS 714 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=304270 $Y=176390 $D=2
M30 714 VSS 4307 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=304270 $Y=328100 $D=2
M31 VSS 4304 4305 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=304720 $Y=177840 $D=2
M32 VSS 4306 4307 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=304720 $Y=326470 $D=2
M33 4304 4305 VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=305860 $Y=177840 $D=2
M34 4306 4307 VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=305860 $Y=326470 $D=2
M35 4304 VSS 713 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=306310 $Y=176390 $D=2
M36 713 VSS 4306 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=306310 $Y=328100 $D=2
M37 4747 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=418270 $Y=176390 $D=2
M38 614 VSS 4749 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=193100 $D=2
M39 4751 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=194390 $D=2
M40 614 VSS 4753 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=211100 $D=2
M41 4755 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=212390 $D=2
M42 614 VSS 4757 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=229100 $D=2
M43 4759 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=230390 $D=2
M44 614 VSS 4761 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=247100 $D=2
M45 4763 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=248390 $D=2
M46 614 VSS 4765 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=265100 $D=2
M47 4767 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=266390 $D=2
M48 614 VSS 4769 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=283100 $D=2
M49 4771 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=284390 $D=2
M50 614 VSS 4773 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=301100 $D=2
M51 4775 VSS 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=302390 $D=2
M52 614 804 4777 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=418270 $Y=319100 $D=2
M53 4743 804 614 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=418270 $Y=320390 $D=2
M54 614 804 4745 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=418270 $Y=328100 $D=2
M55 VSS VDD 4747 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=177840 $D=2
M56 VSS VDD 4749 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=191470 $D=2
M57 VSS VDD 4751 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=195840 $D=2
M58 VSS VDD 4753 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=209470 $D=2
M59 VSS VDD 4755 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=213840 $D=2
M60 VSS VDD 4757 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=227470 $D=2
M61 VSS VDD 4759 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=231840 $D=2
M62 VSS VDD 4761 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=245470 $D=2
M63 VSS VDD 4763 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=249840 $D=2
M64 VSS VDD 4765 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=263470 $D=2
M65 VSS VDD 4767 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=267840 $D=2
M66 VSS VDD 4769 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=281470 $D=2
M67 VSS VDD 4771 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=285840 $D=2
M68 VSS VDD 4773 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=299470 $D=2
M69 VSS VDD 4775 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=303840 $D=2
M70 VSS VDD 4777 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=317470 $D=2
M71 VSS VDD 4743 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=321840 $D=2
M72 VSS VDD 4745 VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.84565e-14 AS=1.18957e-13 PD=-7.88406e-08 PS=9.41159e-07 NRD=0.0204504 NRS=0.131808 m=1 nf=1 $X=418720 $Y=326470 $D=2
M73 4748 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=177840 $D=2
M74 4750 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=191470 $D=2
M75 4752 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=195840 $D=2
M76 4754 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=209470 $D=2
M77 4756 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=213840 $D=2
M78 4758 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=227470 $D=2
M79 4760 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=231840 $D=2
M80 4762 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=245470 $D=2
M81 4764 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=249840 $D=2
M82 4766 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=263470 $D=2
M83 4768 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=267840 $D=2
M84 4770 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=281470 $D=2
M85 4772 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=285840 $D=2
M86 4774 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=299470 $D=2
M87 4776 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=303840 $D=2
M88 4778 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=317470 $D=2
M89 4744 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=321840 $D=2
M90 4746 VSS VSS VSS nfet_05v0 L=6e-07 W=9.5e-07 AD=1.18957e-13 AS=1.84565e-14 PD=9.41159e-07 PS=-7.88406e-08 NRD=0.131808 NRS=0.0204504 m=1 nf=1 $X=419860 $Y=326470 $D=2
M91 606 614 VSS VSS nfet_05v0 L=6e-07 W=2.76e-06 AD=7.176e-13 AS=1.2144e-12 PD=3.8e-06 PS=7.28e-06 NRD=0.376812 NRS=0.637681 m=1 nf=2 $X=418770 $Y=94540 $D=2
M92 607 606 VSS VSS nfet_05v0 L=6e-07 W=1.7e-05 AD=4.42e-12 AS=7.48e-12 PD=1.804e-05 PS=3.576e-05 NRD=0.0611765 NRS=0.103529 m=1 nf=2 $X=418790 $Y=79115 $D=2
M93 613 VDD VSS VSS nfet_05v0 L=6e-07 W=1.14e-06 AD=2.964e-13 AS=5.016e-13 PD=2.18e-06 PS=4.04e-06 NRD=0.912281 NRS=1.54386 m=1 nf=2 $X=419015 $Y=110805 $D=2
M94 4748 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.81613e-13 AS=2.82e-13 PD=1.84258e-06 PS=2.14e-06 NRD=0.782258 NRS=0.783333 m=1 nf=1 $X=420310 $Y=176390 $D=2
M95 615 VSS 4750 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=193100 $D=2
M96 4752 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=194390 $D=2
M97 615 VSS 4754 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=211100 $D=2
M98 4756 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=212390 $D=2
M99 615 VSS 4758 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=229100 $D=2
M100 4760 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=230390 $D=2
M101 615 VSS 4762 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=247100 $D=2
M102 4764 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=248390 $D=2
M103 615 VSS 4766 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=265100 $D=2
M104 4768 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=266390 $D=2
M105 615 VSS 4770 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=283100 $D=2
M106 4772 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=284390 $D=2
M107 615 VSS 4774 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=301100 $D=2
M108 4776 VSS 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=302390 $D=2
M109 615 804 4778 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=-2.739e-13 AS=1.416e-13 PD=-1.70545e-06 PS=8.14545e-07 NRD=-0.760833 NRS=0.393333 m=1 nf=1 $X=420310 $Y=319100 $D=2
M110 4744 804 615 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=1.416e-13 AS=-2.739e-13 PD=8.14545e-07 PS=-1.70545e-06 NRD=0.393333 NRS=-0.760833 m=1 nf=1 $X=420310 $Y=320390 $D=2
M111 615 804 4746 VSS nfet_05v0 L=7.7e-07 W=6e-07 AD=2.82e-13 AS=2.81613e-13 PD=2.14e-06 PS=1.84258e-06 NRD=0.783333 NRS=0.782258 m=1 nf=1 $X=420310 $Y=328100 $D=2
M112 VDD 4249 4251 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=179690 $D=8
M113 VDD 4856 4855 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=180970 $D=8
M114 VDD 4864 4863 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=215690 $D=8
M115 VDD 4920 4919 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=216970 $D=8
M116 VDD 4928 4927 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=251690 $D=8
M117 VDD 4984 4983 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=252970 $D=8
M118 VDD 4992 4991 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=287690 $D=8
M119 VDD 5048 5047 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=288970 $D=8
M120 VDD 5056 5055 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=323690 $D=8
M121 VDD 4337 4339 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=12840 $Y=324970 $D=8
M122 4249 4251 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=179690 $D=8
M123 4856 4855 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=180970 $D=8
M124 4864 4863 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=215690 $D=8
M125 4920 4919 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=216970 $D=8
M126 4928 4927 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=251690 $D=8
M127 4984 4983 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=252970 $D=8
M128 4992 4991 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=287690 $D=8
M129 5048 5047 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=288970 $D=8
M130 5056 5055 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=323690 $D=8
M131 4337 4339 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=13980 $Y=324970 $D=8
M132 4616 4097 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=13620 $Y=160970 $D=8
M133 4617 4097 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=13620 $Y=164845 $D=8
M134 4779 4571 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=13835 $Y=112830 $D=8
M135 VDD 4245 4247 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=179690 $D=8
M136 VDD 4858 4857 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=180970 $D=8
M137 VDD 4866 4865 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=215690 $D=8
M138 VDD 4922 4921 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=216970 $D=8
M139 VDD 4930 4929 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=251690 $D=8
M140 VDD 4986 4985 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=252970 $D=8
M141 VDD 4994 4993 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=287690 $D=8
M142 VDD 5050 5049 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=288970 $D=8
M143 VDD 5058 5057 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=323690 $D=8
M144 VDD 4333 4335 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=15840 $Y=324970 $D=8
M145 4245 4247 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=179690 $D=8
M146 4858 4857 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=180970 $D=8
M147 4866 4865 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=215690 $D=8
M148 4922 4921 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=216970 $D=8
M149 4930 4929 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=251690 $D=8
M150 4986 4985 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=252970 $D=8
M151 4994 4993 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=287690 $D=8
M152 5050 5049 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=288970 $D=8
M153 5058 5057 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=323690 $D=8
M154 4333 4335 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=16980 $Y=324970 $D=8
M155 4780 4570 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=16365 $Y=112830 $D=8
M156 4619 4097 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=16720 $Y=160970 $D=8
M157 4618 4097 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=16720 $Y=164845 $D=8
M158 VDD 4241 4243 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=179690 $D=8
M159 VDD 4860 4859 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=180970 $D=8
M160 VDD 4868 4867 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=215690 $D=8
M161 VDD 4924 4923 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=216970 $D=8
M162 VDD 4932 4931 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=251690 $D=8
M163 VDD 4988 4987 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=252970 $D=8
M164 VDD 4996 4995 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=287690 $D=8
M165 VDD 5052 5051 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=288970 $D=8
M166 VDD 5060 5059 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=323690 $D=8
M167 VDD 4329 4331 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=18840 $Y=324970 $D=8
M168 4241 4243 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=179690 $D=8
M169 4860 4859 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=180970 $D=8
M170 4868 4867 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=215690 $D=8
M171 4924 4923 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=216970 $D=8
M172 4932 4931 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=251690 $D=8
M173 4988 4987 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=252970 $D=8
M174 4996 4995 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=287690 $D=8
M175 5052 5051 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=288970 $D=8
M176 5060 5059 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=323690 $D=8
M177 4329 4331 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=19980 $Y=324970 $D=8
M178 4620 4097 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=19815 $Y=160970 $D=8
M179 4621 4097 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=19815 $Y=164845 $D=8
M180 4781 4569 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=20030 $Y=112830 $D=8
M181 VDD 4237 4239 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=179690 $D=8
M182 VDD 4862 4861 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=180970 $D=8
M183 VDD 4870 4869 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=215690 $D=8
M184 VDD 4926 4925 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=216970 $D=8
M185 VDD 4934 4933 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=251690 $D=8
M186 VDD 4990 4989 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=252970 $D=8
M187 VDD 4998 4997 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=287690 $D=8
M188 VDD 5054 5053 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=288970 $D=8
M189 VDD 5062 5061 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=323690 $D=8
M190 VDD 4325 4327 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=21840 $Y=324970 $D=8
M191 4237 4239 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=179690 $D=8
M192 4862 4861 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=180970 $D=8
M193 4870 4869 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=215690 $D=8
M194 4926 4925 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=216970 $D=8
M195 4934 4933 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=251690 $D=8
M196 4990 4989 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=252970 $D=8
M197 4998 4997 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=287690 $D=8
M198 5054 5053 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=288970 $D=8
M199 5062 5061 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=323690 $D=8
M200 4325 4327 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=22980 $Y=324970 $D=8
M201 4782 4568 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=22560 $Y=112830 $D=8
M202 4623 4097 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=22915 $Y=160970 $D=8
M203 4622 4097 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=22915 $Y=164845 $D=8
M204 VDD 4177 4179 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=179690 $D=8
M205 VDD 4840 4839 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=180970 $D=8
M206 VDD 4848 4847 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=215690 $D=8
M207 VDD 4904 4903 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=216970 $D=8
M208 VDD 4912 4911 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=251690 $D=8
M209 VDD 4968 4967 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=252970 $D=8
M210 VDD 4976 4975 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=287690 $D=8
M211 VDD 5032 5031 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=288970 $D=8
M212 VDD 5040 5039 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=323690 $D=8
M213 VDD 4321 4323 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=24840 $Y=324970 $D=8
M214 4177 4179 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=179690 $D=8
M215 4840 4839 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=180970 $D=8
M216 4848 4847 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=215690 $D=8
M217 4904 4903 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=216970 $D=8
M218 4912 4911 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=251690 $D=8
M219 4968 4967 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=252970 $D=8
M220 4976 4975 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=287690 $D=8
M221 5032 5031 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=288970 $D=8
M222 5040 5039 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=323690 $D=8
M223 4321 4323 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=25980 $Y=324970 $D=8
M224 4624 4097 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=26005 $Y=160970 $D=8
M225 4625 4097 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=26005 $Y=164845 $D=8
M226 4783 4567 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=26220 $Y=112830 $D=8
M227 VDD 4173 4175 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=179690 $D=8
M228 VDD 4842 4841 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=180970 $D=8
M229 VDD 4850 4849 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=215690 $D=8
M230 VDD 4906 4905 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=216970 $D=8
M231 VDD 4914 4913 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=251690 $D=8
M232 VDD 4970 4969 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=252970 $D=8
M233 VDD 4978 4977 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=287690 $D=8
M234 VDD 5034 5033 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=288970 $D=8
M235 VDD 5042 5041 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=323690 $D=8
M236 VDD 4317 4319 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=27840 $Y=324970 $D=8
M237 4173 4175 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=179690 $D=8
M238 4842 4841 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=180970 $D=8
M239 4850 4849 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=215690 $D=8
M240 4906 4905 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=216970 $D=8
M241 4914 4913 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=251690 $D=8
M242 4970 4969 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=252970 $D=8
M243 4978 4977 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=287690 $D=8
M244 5034 5033 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=288970 $D=8
M245 5042 5041 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=323690 $D=8
M246 4317 4319 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=28980 $Y=324970 $D=8
M247 4784 4566 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=28750 $Y=112830 $D=8
M248 4627 4097 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=29105 $Y=160970 $D=8
M249 4626 4097 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=29105 $Y=164845 $D=8
M250 VDD 4185 4187 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=179690 $D=8
M251 VDD 4844 4843 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=180970 $D=8
M252 VDD 4852 4851 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=215690 $D=8
M253 VDD 4908 4907 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=216970 $D=8
M254 VDD 4916 4915 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=251690 $D=8
M255 VDD 4972 4971 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=252970 $D=8
M256 VDD 4980 4979 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=287690 $D=8
M257 VDD 5036 5035 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=288970 $D=8
M258 VDD 5044 5043 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=323690 $D=8
M259 VDD 4313 4315 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=30840 $Y=324970 $D=8
M260 4185 4187 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=179690 $D=8
M261 4844 4843 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=180970 $D=8
M262 4852 4851 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=215690 $D=8
M263 4908 4907 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=216970 $D=8
M264 4916 4915 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=251690 $D=8
M265 4972 4971 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=252970 $D=8
M266 4980 4979 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=287690 $D=8
M267 5036 5035 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=288970 $D=8
M268 5044 5043 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=323690 $D=8
M269 4313 4315 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=31980 $Y=324970 $D=8
M270 4628 4097 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=32200 $Y=160970 $D=8
M271 4629 4097 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=32200 $Y=164845 $D=8
M272 4785 4565 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=32415 $Y=112830 $D=8
M273 VDD 4181 4183 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=179690 $D=8
M274 VDD 4846 4845 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=180970 $D=8
M275 VDD 4854 4853 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=215690 $D=8
M276 VDD 4910 4909 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=216970 $D=8
M277 VDD 4918 4917 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=251690 $D=8
M278 VDD 4974 4973 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=252970 $D=8
M279 VDD 4982 4981 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=287690 $D=8
M280 VDD 5038 5037 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=288970 $D=8
M281 VDD 5046 5045 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=323690 $D=8
M282 VDD 4309 4311 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=33840 $Y=324970 $D=8
M283 4181 4183 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=179690 $D=8
M284 4846 4845 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=180970 $D=8
M285 4854 4853 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=215690 $D=8
M286 4910 4909 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=216970 $D=8
M287 4918 4917 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=251690 $D=8
M288 4974 4973 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=252970 $D=8
M289 4982 4981 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=287690 $D=8
M290 5038 5037 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=288970 $D=8
M291 5046 5045 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=323690 $D=8
M292 4309 4311 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=34980 $Y=324970 $D=8
M293 4735 4564 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=34945 $Y=112830 $D=8
M294 881 4097 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=35120 $Y=160970 $D=8
M295 882 4097 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=35120 $Y=164845 $D=8
M296 893 891 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=38575 $Y=160970 $D=8
M297 894 891 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=38575 $Y=164845 $D=8
M298 VDD 4369 4371 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=179690 $D=8
M299 VDD 4829 4830 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=180970 $D=8
M300 VDD 4837 4838 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=215690 $D=8
M301 VDD 4893 4894 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=216970 $D=8
M302 VDD 4901 4902 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=251690 $D=8
M303 VDD 4957 4958 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=252970 $D=8
M304 VDD 4965 4966 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=287690 $D=8
M305 VDD 5021 5022 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=288970 $D=8
M306 VDD 5029 5030 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=323690 $D=8
M307 VDD 4401 4403 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=39840 $Y=324970 $D=8
M308 4739 4571 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=38620 $Y=112830 $D=8
M309 4369 4371 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=179690 $D=8
M310 4829 4830 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=180970 $D=8
M311 4837 4838 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=215690 $D=8
M312 4893 4894 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=216970 $D=8
M313 4901 4902 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=251690 $D=8
M314 4957 4958 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=252970 $D=8
M315 4965 4966 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=287690 $D=8
M316 5021 5022 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=288970 $D=8
M317 5029 5030 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=323690 $D=8
M318 4401 4403 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=40980 $Y=324970 $D=8
M319 5325 4570 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=41145 $Y=112830 $D=8
M320 4684 891 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=41500 $Y=160970 $D=8
M321 4685 891 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=41500 $Y=164845 $D=8
M322 VDD 4365 4367 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=179690 $D=8
M323 VDD 4827 4828 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=180970 $D=8
M324 VDD 4835 4836 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=215690 $D=8
M325 VDD 4891 4892 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=216970 $D=8
M326 VDD 4899 4900 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=251690 $D=8
M327 VDD 4955 4956 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=252970 $D=8
M328 VDD 4963 4964 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=287690 $D=8
M329 VDD 5019 5020 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=288970 $D=8
M330 VDD 5027 5028 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=323690 $D=8
M331 VDD 4397 4399 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=42840 $Y=324970 $D=8
M332 4365 4367 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=179690 $D=8
M333 4827 4828 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=180970 $D=8
M334 4835 4836 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=215690 $D=8
M335 4891 4892 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=216970 $D=8
M336 4899 4900 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=251690 $D=8
M337 4955 4956 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=252970 $D=8
M338 4963 4964 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=287690 $D=8
M339 5019 5020 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=288970 $D=8
M340 5027 5028 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=323690 $D=8
M341 4397 4399 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=43980 $Y=324970 $D=8
M342 4683 891 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=44595 $Y=160970 $D=8
M343 4682 891 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=44595 $Y=164845 $D=8
M344 VDD 4361 4363 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=179690 $D=8
M345 VDD 4825 4826 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=180970 $D=8
M346 VDD 4833 4834 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=215690 $D=8
M347 VDD 4889 4890 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=216970 $D=8
M348 VDD 4897 4898 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=251690 $D=8
M349 VDD 4953 4954 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=252970 $D=8
M350 VDD 4961 4962 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=287690 $D=8
M351 VDD 5017 5018 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=288970 $D=8
M352 VDD 5025 5026 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=323690 $D=8
M353 VDD 4393 4395 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=45840 $Y=324970 $D=8
M354 5324 4569 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=44810 $Y=112830 $D=8
M355 4361 4363 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=179690 $D=8
M356 4825 4826 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=180970 $D=8
M357 4833 4834 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=215690 $D=8
M358 4889 4890 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=216970 $D=8
M359 4897 4898 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=251690 $D=8
M360 4953 4954 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=252970 $D=8
M361 4961 4962 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=287690 $D=8
M362 5017 5018 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=288970 $D=8
M363 5025 5026 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=323690 $D=8
M364 4393 4395 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=46980 $Y=324970 $D=8
M365 5323 4568 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=47340 $Y=112830 $D=8
M366 4680 891 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=47695 $Y=160970 $D=8
M367 4681 891 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=47695 $Y=164845 $D=8
M368 VDD 4357 4359 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=179690 $D=8
M369 VDD 4823 4824 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=180970 $D=8
M370 VDD 4831 4832 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=215690 $D=8
M371 VDD 4887 4888 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=216970 $D=8
M372 VDD 4895 4896 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=251690 $D=8
M373 VDD 4951 4952 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=252970 $D=8
M374 VDD 4959 4960 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=287690 $D=8
M375 VDD 5015 5016 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=288970 $D=8
M376 VDD 5023 5024 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=323690 $D=8
M377 VDD 4389 4391 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=48840 $Y=324970 $D=8
M378 4357 4359 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=179690 $D=8
M379 4823 4824 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=180970 $D=8
M380 4831 4832 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=215690 $D=8
M381 4887 4888 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=216970 $D=8
M382 4895 4896 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=251690 $D=8
M383 4951 4952 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=252970 $D=8
M384 4959 4960 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=287690 $D=8
M385 5015 5016 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=288970 $D=8
M386 5023 5024 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=323690 $D=8
M387 4389 4391 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=49980 $Y=324970 $D=8
M388 VDD 4353 4355 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=179690 $D=8
M389 VDD 4813 4814 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=180970 $D=8
M390 VDD 4821 4822 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=215690 $D=8
M391 VDD 4877 4878 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=216970 $D=8
M392 VDD 4885 4886 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=251690 $D=8
M393 VDD 4941 4942 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=252970 $D=8
M394 VDD 4949 4950 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=287690 $D=8
M395 VDD 5005 5006 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=288970 $D=8
M396 VDD 5013 5014 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=323690 $D=8
M397 VDD 4385 4387 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=51840 $Y=324970 $D=8
M398 4679 891 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=50785 $Y=160970 $D=8
M399 4678 891 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=50785 $Y=164845 $D=8
M400 5322 4567 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=51000 $Y=112830 $D=8
M401 4353 4355 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=179690 $D=8
M402 4813 4814 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=180970 $D=8
M403 4821 4822 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=215690 $D=8
M404 4877 4878 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=216970 $D=8
M405 4885 4886 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=251690 $D=8
M406 4941 4942 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=252970 $D=8
M407 4949 4950 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=287690 $D=8
M408 5005 5006 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=288970 $D=8
M409 5013 5014 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=323690 $D=8
M410 4385 4387 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=52980 $Y=324970 $D=8
M411 5321 4566 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=53530 $Y=112830 $D=8
M412 VDD 4349 4351 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=179690 $D=8
M413 VDD 4811 4812 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=180970 $D=8
M414 VDD 4819 4820 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=215690 $D=8
M415 VDD 4875 4876 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=216970 $D=8
M416 VDD 4883 4884 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=251690 $D=8
M417 VDD 4939 4940 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=252970 $D=8
M418 VDD 4947 4948 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=287690 $D=8
M419 VDD 5003 5004 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=288970 $D=8
M420 VDD 5011 5012 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=323690 $D=8
M421 VDD 4381 4383 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=54840 $Y=324970 $D=8
M422 4676 891 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=53885 $Y=160970 $D=8
M423 4677 891 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=53885 $Y=164845 $D=8
M424 4349 4351 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=179690 $D=8
M425 4811 4812 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=180970 $D=8
M426 4819 4820 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=215690 $D=8
M427 4875 4876 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=216970 $D=8
M428 4883 4884 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=251690 $D=8
M429 4939 4940 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=252970 $D=8
M430 4947 4948 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=287690 $D=8
M431 5003 5004 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=288970 $D=8
M432 5011 5012 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=323690 $D=8
M433 4381 4383 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=55980 $Y=324970 $D=8
M434 VDD 4345 4347 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=179690 $D=8
M435 VDD 4809 4810 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=180970 $D=8
M436 VDD 4817 4818 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=215690 $D=8
M437 VDD 4873 4874 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=216970 $D=8
M438 VDD 4881 4882 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=251690 $D=8
M439 VDD 4937 4938 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=252970 $D=8
M440 VDD 4945 4946 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=287690 $D=8
M441 VDD 5001 5002 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=288970 $D=8
M442 VDD 5009 5010 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=323690 $D=8
M443 VDD 4377 4379 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=57840 $Y=324970 $D=8
M444 4675 891 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=56980 $Y=160970 $D=8
M445 4674 891 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=56980 $Y=164845 $D=8
M446 5320 4565 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=57195 $Y=112830 $D=8
M447 4345 4347 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=179690 $D=8
M448 4809 4810 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=180970 $D=8
M449 4817 4818 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=215690 $D=8
M450 4873 4874 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=216970 $D=8
M451 4881 4882 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=251690 $D=8
M452 4937 4938 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=252970 $D=8
M453 4945 4946 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=287690 $D=8
M454 5001 5002 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=288970 $D=8
M455 5009 5010 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=323690 $D=8
M456 4377 4379 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=58980 $Y=324970 $D=8
M457 VDD 4341 4343 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=179690 $D=8
M458 VDD 4807 4808 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=180970 $D=8
M459 VDD 4815 4816 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=215690 $D=8
M460 VDD 4871 4872 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=216970 $D=8
M461 VDD 4879 4880 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=251690 $D=8
M462 VDD 4935 4936 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=252970 $D=8
M463 VDD 4943 4944 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=287690 $D=8
M464 VDD 4999 5000 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=288970 $D=8
M465 VDD 5007 5008 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=323690 $D=8
M466 VDD 4373 4375 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=60840 $Y=324970 $D=8
M467 5319 4564 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=59725 $Y=112830 $D=8
M468 4672 891 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=60080 $Y=160970 $D=8
M469 4673 891 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=60080 $Y=164845 $D=8
M470 4341 4343 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=179690 $D=8
M471 4807 4808 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=180970 $D=8
M472 4815 4816 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=215690 $D=8
M473 4871 4872 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=216970 $D=8
M474 4879 4880 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=251690 $D=8
M475 4935 4936 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=252970 $D=8
M476 4943 4944 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=287690 $D=8
M477 4999 5000 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=288970 $D=8
M478 5007 5008 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=323690 $D=8
M479 4373 4375 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=61980 $Y=324970 $D=8
M480 VDD 4265 4267 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=179690 $D=8
M481 VDD 5112 5111 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=180970 $D=8
M482 VDD 5120 5119 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=215690 $D=8
M483 VDD 5176 5175 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=216970 $D=8
M484 VDD 5184 5183 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=251690 $D=8
M485 VDD 5240 5239 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=252970 $D=8
M486 VDD 5248 5247 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=287690 $D=8
M487 VDD 5304 5303 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=288970 $D=8
M488 VDD 5312 5311 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=323690 $D=8
M489 VDD 4433 4435 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=66840 $Y=324970 $D=8
M490 4265 4267 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=179690 $D=8
M491 5112 5111 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=180970 $D=8
M492 5120 5119 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=215690 $D=8
M493 5176 5175 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=216970 $D=8
M494 5184 5183 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=251690 $D=8
M495 5240 5239 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=252970 $D=8
M496 5248 5247 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=287690 $D=8
M497 5304 5303 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=288970 $D=8
M498 5312 5311 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=323690 $D=8
M499 4433 4435 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=67980 $Y=324970 $D=8
M500 4630 4098 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=67620 $Y=160970 $D=8
M501 4631 4098 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=67620 $Y=164845 $D=8
M502 4786 4571 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=67835 $Y=112830 $D=8
M503 VDD 4261 4263 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=179690 $D=8
M504 VDD 5114 5113 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=180970 $D=8
M505 VDD 5122 5121 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=215690 $D=8
M506 VDD 5178 5177 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=216970 $D=8
M507 VDD 5186 5185 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=251690 $D=8
M508 VDD 5242 5241 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=252970 $D=8
M509 VDD 5250 5249 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=287690 $D=8
M510 VDD 5306 5305 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=288970 $D=8
M511 VDD 5314 5313 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=323690 $D=8
M512 VDD 4429 4431 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=69840 $Y=324970 $D=8
M513 4261 4263 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=179690 $D=8
M514 5114 5113 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=180970 $D=8
M515 5122 5121 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=215690 $D=8
M516 5178 5177 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=216970 $D=8
M517 5186 5185 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=251690 $D=8
M518 5242 5241 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=252970 $D=8
M519 5250 5249 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=287690 $D=8
M520 5306 5305 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=288970 $D=8
M521 5314 5313 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=323690 $D=8
M522 4429 4431 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=70980 $Y=324970 $D=8
M523 4787 4570 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=70365 $Y=112830 $D=8
M524 4633 4098 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=70720 $Y=160970 $D=8
M525 4632 4098 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=70720 $Y=164845 $D=8
M526 VDD 4257 4259 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=179690 $D=8
M527 VDD 5116 5115 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=180970 $D=8
M528 VDD 5124 5123 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=215690 $D=8
M529 VDD 5180 5179 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=216970 $D=8
M530 VDD 5188 5187 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=251690 $D=8
M531 VDD 5244 5243 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=252970 $D=8
M532 VDD 5252 5251 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=287690 $D=8
M533 VDD 5308 5307 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=288970 $D=8
M534 VDD 5316 5315 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=323690 $D=8
M535 VDD 4425 4427 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=72840 $Y=324970 $D=8
M536 4257 4259 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=179690 $D=8
M537 5116 5115 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=180970 $D=8
M538 5124 5123 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=215690 $D=8
M539 5180 5179 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=216970 $D=8
M540 5188 5187 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=251690 $D=8
M541 5244 5243 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=252970 $D=8
M542 5252 5251 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=287690 $D=8
M543 5308 5307 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=288970 $D=8
M544 5316 5315 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=323690 $D=8
M545 4425 4427 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=73980 $Y=324970 $D=8
M546 4634 4098 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=73815 $Y=160970 $D=8
M547 4635 4098 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=73815 $Y=164845 $D=8
M548 4788 4569 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=74030 $Y=112830 $D=8
M549 VDD 4253 4255 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=179690 $D=8
M550 VDD 5118 5117 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=180970 $D=8
M551 VDD 5126 5125 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=215690 $D=8
M552 VDD 5182 5181 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=216970 $D=8
M553 VDD 5190 5189 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=251690 $D=8
M554 VDD 5246 5245 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=252970 $D=8
M555 VDD 5254 5253 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=287690 $D=8
M556 VDD 5310 5309 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=288970 $D=8
M557 VDD 5318 5317 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=323690 $D=8
M558 VDD 4421 4423 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=75840 $Y=324970 $D=8
M559 4253 4255 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=179690 $D=8
M560 5118 5117 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=180970 $D=8
M561 5126 5125 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=215690 $D=8
M562 5182 5181 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=216970 $D=8
M563 5190 5189 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=251690 $D=8
M564 5246 5245 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=252970 $D=8
M565 5254 5253 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=287690 $D=8
M566 5310 5309 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=288970 $D=8
M567 5318 5317 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=323690 $D=8
M568 4421 4423 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=76980 $Y=324970 $D=8
M569 4789 4568 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=76560 $Y=112830 $D=8
M570 4637 4098 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=76915 $Y=160970 $D=8
M571 4636 4098 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=76915 $Y=164845 $D=8
M572 VDD 4193 4195 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=179690 $D=8
M573 VDD 5096 5095 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=180970 $D=8
M574 VDD 5104 5103 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=215690 $D=8
M575 VDD 5160 5159 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=216970 $D=8
M576 VDD 5168 5167 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=251690 $D=8
M577 VDD 5224 5223 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=252970 $D=8
M578 VDD 5232 5231 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=287690 $D=8
M579 VDD 5288 5287 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=288970 $D=8
M580 VDD 5296 5295 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=323690 $D=8
M581 VDD 4417 4419 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=78840 $Y=324970 $D=8
M582 4193 4195 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=179690 $D=8
M583 5096 5095 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=180970 $D=8
M584 5104 5103 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=215690 $D=8
M585 5160 5159 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=216970 $D=8
M586 5168 5167 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=251690 $D=8
M587 5224 5223 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=252970 $D=8
M588 5232 5231 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=287690 $D=8
M589 5288 5287 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=288970 $D=8
M590 5296 5295 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=323690 $D=8
M591 4417 4419 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=79980 $Y=324970 $D=8
M592 4638 4098 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=80005 $Y=160970 $D=8
M593 4639 4098 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=80005 $Y=164845 $D=8
M594 4790 4567 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=80220 $Y=112830 $D=8
M595 VDD 4189 4191 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=179690 $D=8
M596 VDD 5098 5097 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=180970 $D=8
M597 VDD 5106 5105 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=215690 $D=8
M598 VDD 5162 5161 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=216970 $D=8
M599 VDD 5170 5169 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=251690 $D=8
M600 VDD 5226 5225 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=252970 $D=8
M601 VDD 5234 5233 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=287690 $D=8
M602 VDD 5290 5289 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=288970 $D=8
M603 VDD 5298 5297 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=323690 $D=8
M604 VDD 4413 4415 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=81840 $Y=324970 $D=8
M605 4189 4191 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=179690 $D=8
M606 5098 5097 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=180970 $D=8
M607 5106 5105 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=215690 $D=8
M608 5162 5161 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=216970 $D=8
M609 5170 5169 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=251690 $D=8
M610 5226 5225 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=252970 $D=8
M611 5234 5233 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=287690 $D=8
M612 5290 5289 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=288970 $D=8
M613 5298 5297 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=323690 $D=8
M614 4413 4415 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=82980 $Y=324970 $D=8
M615 4791 4566 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=82750 $Y=112830 $D=8
M616 4641 4098 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=83105 $Y=160970 $D=8
M617 4640 4098 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=83105 $Y=164845 $D=8
M618 VDD 4201 4203 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=179690 $D=8
M619 VDD 5100 5099 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=180970 $D=8
M620 VDD 5108 5107 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=215690 $D=8
M621 VDD 5164 5163 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=216970 $D=8
M622 VDD 5172 5171 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=251690 $D=8
M623 VDD 5228 5227 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=252970 $D=8
M624 VDD 5236 5235 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=287690 $D=8
M625 VDD 5292 5291 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=288970 $D=8
M626 VDD 5300 5299 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=323690 $D=8
M627 VDD 4409 4411 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=84840 $Y=324970 $D=8
M628 4201 4203 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=179690 $D=8
M629 5100 5099 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=180970 $D=8
M630 5108 5107 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=215690 $D=8
M631 5164 5163 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=216970 $D=8
M632 5172 5171 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=251690 $D=8
M633 5228 5227 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=252970 $D=8
M634 5236 5235 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=287690 $D=8
M635 5292 5291 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=288970 $D=8
M636 5300 5299 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=323690 $D=8
M637 4409 4411 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=85980 $Y=324970 $D=8
M638 4642 4098 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=86200 $Y=160970 $D=8
M639 4643 4098 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=86200 $Y=164845 $D=8
M640 4792 4565 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=86415 $Y=112830 $D=8
M641 VDD 4197 4199 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=179690 $D=8
M642 VDD 5102 5101 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=180970 $D=8
M643 VDD 5110 5109 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=215690 $D=8
M644 VDD 5166 5165 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=216970 $D=8
M645 VDD 5174 5173 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=251690 $D=8
M646 VDD 5230 5229 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=252970 $D=8
M647 VDD 5238 5237 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=287690 $D=8
M648 VDD 5294 5293 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=288970 $D=8
M649 VDD 5302 5301 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=323690 $D=8
M650 VDD 4405 4407 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=87840 $Y=324970 $D=8
M651 4197 4199 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=179690 $D=8
M652 5102 5101 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=180970 $D=8
M653 5110 5109 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=215690 $D=8
M654 5166 5165 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=216970 $D=8
M655 5174 5173 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=251690 $D=8
M656 5230 5229 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=252970 $D=8
M657 5238 5237 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=287690 $D=8
M658 5294 5293 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=288970 $D=8
M659 5302 5301 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=323690 $D=8
M660 4405 4407 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=88980 $Y=324970 $D=8
M661 4736 4564 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=88945 $Y=112830 $D=8
M662 883 4098 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=89120 $Y=160970 $D=8
M663 884 4098 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=89120 $Y=164845 $D=8
M664 896 895 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=92575 $Y=160970 $D=8
M665 897 895 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=92575 $Y=164845 $D=8
M666 VDD 4465 4467 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=179690 $D=8
M667 VDD 5085 5086 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=180970 $D=8
M668 VDD 5093 5094 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=215690 $D=8
M669 VDD 5149 5150 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=216970 $D=8
M670 VDD 5157 5158 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=251690 $D=8
M671 VDD 5213 5214 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=252970 $D=8
M672 VDD 5221 5222 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=287690 $D=8
M673 VDD 5277 5278 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=288970 $D=8
M674 VDD 5285 5286 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=323690 $D=8
M675 VDD 4497 4499 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=93840 $Y=324970 $D=8
M676 4740 4571 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=92620 $Y=112830 $D=8
M677 4465 4467 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=179690 $D=8
M678 5085 5086 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=180970 $D=8
M679 5093 5094 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=215690 $D=8
M680 5149 5150 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=216970 $D=8
M681 5157 5158 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=251690 $D=8
M682 5213 5214 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=252970 $D=8
M683 5221 5222 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=287690 $D=8
M684 5277 5278 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=288970 $D=8
M685 5285 5286 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=323690 $D=8
M686 4497 4499 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=94980 $Y=324970 $D=8
M687 5332 4570 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=95145 $Y=112830 $D=8
M688 4698 895 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=95500 $Y=160970 $D=8
M689 4699 895 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=95500 $Y=164845 $D=8
M690 VDD 4461 4463 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=179690 $D=8
M691 VDD 5083 5084 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=180970 $D=8
M692 VDD 5091 5092 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=215690 $D=8
M693 VDD 5147 5148 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=216970 $D=8
M694 VDD 5155 5156 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=251690 $D=8
M695 VDD 5211 5212 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=252970 $D=8
M696 VDD 5219 5220 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=287690 $D=8
M697 VDD 5275 5276 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=288970 $D=8
M698 VDD 5283 5284 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=323690 $D=8
M699 VDD 4493 4495 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=96840 $Y=324970 $D=8
M700 4461 4463 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=179690 $D=8
M701 5083 5084 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=180970 $D=8
M702 5091 5092 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=215690 $D=8
M703 5147 5148 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=216970 $D=8
M704 5155 5156 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=251690 $D=8
M705 5211 5212 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=252970 $D=8
M706 5219 5220 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=287690 $D=8
M707 5275 5276 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=288970 $D=8
M708 5283 5284 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=323690 $D=8
M709 4493 4495 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=97980 $Y=324970 $D=8
M710 4697 895 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=98595 $Y=160970 $D=8
M711 4696 895 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=98595 $Y=164845 $D=8
M712 VDD 4457 4459 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=179690 $D=8
M713 VDD 5081 5082 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=180970 $D=8
M714 VDD 5089 5090 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=215690 $D=8
M715 VDD 5145 5146 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=216970 $D=8
M716 VDD 5153 5154 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=251690 $D=8
M717 VDD 5209 5210 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=252970 $D=8
M718 VDD 5217 5218 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=287690 $D=8
M719 VDD 5273 5274 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=288970 $D=8
M720 VDD 5281 5282 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=323690 $D=8
M721 VDD 4489 4491 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=99840 $Y=324970 $D=8
M722 5331 4569 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=98810 $Y=112830 $D=8
M723 4457 4459 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=179690 $D=8
M724 5081 5082 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=180970 $D=8
M725 5089 5090 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=215690 $D=8
M726 5145 5146 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=216970 $D=8
M727 5153 5154 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=251690 $D=8
M728 5209 5210 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=252970 $D=8
M729 5217 5218 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=287690 $D=8
M730 5273 5274 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=288970 $D=8
M731 5281 5282 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=323690 $D=8
M732 4489 4491 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=100980 $Y=324970 $D=8
M733 5330 4568 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=101340 $Y=112830 $D=8
M734 4694 895 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=101695 $Y=160970 $D=8
M735 4695 895 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=101695 $Y=164845 $D=8
M736 VDD 4453 4455 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=179690 $D=8
M737 VDD 5079 5080 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=180970 $D=8
M738 VDD 5087 5088 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=215690 $D=8
M739 VDD 5143 5144 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=216970 $D=8
M740 VDD 5151 5152 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=251690 $D=8
M741 VDD 5207 5208 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=252970 $D=8
M742 VDD 5215 5216 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=287690 $D=8
M743 VDD 5271 5272 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=288970 $D=8
M744 VDD 5279 5280 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=323690 $D=8
M745 VDD 4485 4487 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=102840 $Y=324970 $D=8
M746 4453 4455 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=179690 $D=8
M747 5079 5080 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=180970 $D=8
M748 5087 5088 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=215690 $D=8
M749 5143 5144 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=216970 $D=8
M750 5151 5152 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=251690 $D=8
M751 5207 5208 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=252970 $D=8
M752 5215 5216 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=287690 $D=8
M753 5271 5272 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=288970 $D=8
M754 5279 5280 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=323690 $D=8
M755 4485 4487 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=103980 $Y=324970 $D=8
M756 VDD 4449 4451 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=179690 $D=8
M757 VDD 5069 5070 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=180970 $D=8
M758 VDD 5077 5078 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=215690 $D=8
M759 VDD 5133 5134 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=216970 $D=8
M760 VDD 5141 5142 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=251690 $D=8
M761 VDD 5197 5198 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=252970 $D=8
M762 VDD 5205 5206 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=287690 $D=8
M763 VDD 5261 5262 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=288970 $D=8
M764 VDD 5269 5270 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=323690 $D=8
M765 VDD 4481 4483 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=105840 $Y=324970 $D=8
M766 4693 895 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=104785 $Y=160970 $D=8
M767 4692 895 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=104785 $Y=164845 $D=8
M768 5329 4567 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=105000 $Y=112830 $D=8
M769 4449 4451 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=179690 $D=8
M770 5069 5070 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=180970 $D=8
M771 5077 5078 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=215690 $D=8
M772 5133 5134 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=216970 $D=8
M773 5141 5142 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=251690 $D=8
M774 5197 5198 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=252970 $D=8
M775 5205 5206 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=287690 $D=8
M776 5261 5262 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=288970 $D=8
M777 5269 5270 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=323690 $D=8
M778 4481 4483 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=106980 $Y=324970 $D=8
M779 5328 4566 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=107530 $Y=112830 $D=8
M780 VDD 4445 4447 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=179690 $D=8
M781 VDD 5067 5068 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=180970 $D=8
M782 VDD 5075 5076 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=215690 $D=8
M783 VDD 5131 5132 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=216970 $D=8
M784 VDD 5139 5140 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=251690 $D=8
M785 VDD 5195 5196 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=252970 $D=8
M786 VDD 5203 5204 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=287690 $D=8
M787 VDD 5259 5260 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=288970 $D=8
M788 VDD 5267 5268 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=323690 $D=8
M789 VDD 4477 4479 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=108840 $Y=324970 $D=8
M790 4690 895 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=107885 $Y=160970 $D=8
M791 4691 895 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=107885 $Y=164845 $D=8
M792 4445 4447 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=179690 $D=8
M793 5067 5068 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=180970 $D=8
M794 5075 5076 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=215690 $D=8
M795 5131 5132 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=216970 $D=8
M796 5139 5140 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=251690 $D=8
M797 5195 5196 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=252970 $D=8
M798 5203 5204 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=287690 $D=8
M799 5259 5260 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=288970 $D=8
M800 5267 5268 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=323690 $D=8
M801 4477 4479 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=109980 $Y=324970 $D=8
M802 VDD 4441 4443 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=179690 $D=8
M803 VDD 5065 5066 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=180970 $D=8
M804 VDD 5073 5074 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=215690 $D=8
M805 VDD 5129 5130 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=216970 $D=8
M806 VDD 5137 5138 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=251690 $D=8
M807 VDD 5193 5194 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=252970 $D=8
M808 VDD 5201 5202 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=287690 $D=8
M809 VDD 5257 5258 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=288970 $D=8
M810 VDD 5265 5266 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=323690 $D=8
M811 VDD 4473 4475 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=111840 $Y=324970 $D=8
M812 4689 895 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=110980 $Y=160970 $D=8
M813 4688 895 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=110980 $Y=164845 $D=8
M814 5327 4565 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=111195 $Y=112830 $D=8
M815 4441 4443 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=179690 $D=8
M816 5065 5066 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=180970 $D=8
M817 5073 5074 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=215690 $D=8
M818 5129 5130 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=216970 $D=8
M819 5137 5138 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=251690 $D=8
M820 5193 5194 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=252970 $D=8
M821 5201 5202 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=287690 $D=8
M822 5257 5258 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=288970 $D=8
M823 5265 5266 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=323690 $D=8
M824 4473 4475 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=112980 $Y=324970 $D=8
M825 VDD 4437 4439 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=179690 $D=8
M826 VDD 5063 5064 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=180970 $D=8
M827 VDD 5071 5072 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=215690 $D=8
M828 VDD 5127 5128 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=216970 $D=8
M829 VDD 5135 5136 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=251690 $D=8
M830 VDD 5191 5192 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=252970 $D=8
M831 VDD 5199 5200 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=287690 $D=8
M832 VDD 5255 5256 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=288970 $D=8
M833 VDD 5263 5264 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=323690 $D=8
M834 VDD 4469 4471 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=114840 $Y=324970 $D=8
M835 5326 4564 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=113725 $Y=112830 $D=8
M836 4686 895 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=114080 $Y=160970 $D=8
M837 4687 895 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=114080 $Y=164845 $D=8
M838 4437 4439 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=179690 $D=8
M839 5063 5064 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=180970 $D=8
M840 5071 5072 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=215690 $D=8
M841 5127 5128 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=216970 $D=8
M842 5135 5136 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=251690 $D=8
M843 5191 5192 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=252970 $D=8
M844 5199 5200 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=287690 $D=8
M845 5255 5256 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=288970 $D=8
M846 5263 5264 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=323690 $D=8
M847 4469 4471 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=115980 $Y=324970 $D=8
M848 VDD 4300 4301 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=179690 $D=8
M849 VDD 5349 5350 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=180970 $D=8
M850 VDD 5347 5348 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=188690 $D=8
M851 VDD 5357 5358 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=189970 $D=8
M852 VDD 5355 5356 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=206690 $D=8
M853 VDD 5361 5362 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=207970 $D=8
M854 VDD 5359 5360 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=224690 $D=8
M855 VDD 5365 5366 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=225970 $D=8
M856 VDD 5363 5364 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=242690 $D=8
M857 VDD 5369 5370 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=243970 $D=8
M858 VDD 5367 5368 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=260690 $D=8
M859 VDD 5373 5374 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=261970 $D=8
M860 VDD 5371 5372 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=278690 $D=8
M861 VDD 5377 5378 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=279970 $D=8
M862 VDD 5375 5376 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=296690 $D=8
M863 VDD 5381 5382 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=297970 $D=8
M864 VDD 5379 5380 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=314690 $D=8
M865 VDD 5353 5354 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=315970 $D=8
M866 VDD 5351 5352 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=323690 $D=8
M867 VDD 4302 4303 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=120840 $Y=324970 $D=8
M868 VDD VSS VDD VDD pfet_05v0 L=2.365e-06 W=8.19e-05 AD=0 AS=6.1309e-11 PD=0 PS=0.000217698 NRD=0 NRS=11.8457 m=1 nf=36 $X=10835 $Y=171065 $D=8
M869 4300 4301 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=179690 $D=8
M870 5349 5350 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=180970 $D=8
M871 5347 5348 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=188690 $D=8
M872 5357 5358 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=189970 $D=8
M873 5355 5356 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=206690 $D=8
M874 5361 5362 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=207970 $D=8
M875 5359 5360 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=224690 $D=8
M876 5365 5366 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=225970 $D=8
M877 5363 5364 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=242690 $D=8
M878 5369 5370 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=243970 $D=8
M879 5367 5368 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=260690 $D=8
M880 5373 5374 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=261970 $D=8
M881 5371 5372 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=278690 $D=8
M882 5377 5378 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=279970 $D=8
M883 5375 5376 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=296690 $D=8
M884 5381 5382 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=297970 $D=8
M885 5379 5380 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=314690 $D=8
M886 5353 5354 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=315970 $D=8
M887 5351 5352 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=323690 $D=8
M888 4302 4303 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=121980 $Y=324970 $D=8
M889 VDD VSS VDD VDD pfet_05v0 L=3.94e-06 W=0.000181335 AD=0 AS=1.05339e-10 PD=0 PS=0.000412 NRD=0 NRS=3.48863 m=1 nf=33 $X=146370 $Y=180915 $D=8
M890 4734 1 VDD VDD pfet_05v0 L=5.95e-07 W=2.28e-06 AD=5.985e-13 AS=1.3566e-12 PD=2.805e-06 PS=5.75e-06 NRD=0.115132 NRS=0.260965 m=1 nf=1 $X=233770 $Y=57780 $D=8
M891 617 802 VDD VDD pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=233770 $Y=63100 $D=8
M892 802 CLK 4734 VDD pfet_05v0 L=5.95e-07 W=2.28e-06 AD=1.3566e-12 AS=5.985e-13 PD=5.75e-06 PS=2.805e-06 NRD=0.260965 NRS=0.115132 m=1 nf=1 $X=234890 $Y=57780 $D=8
M893 616 619 VDD VDD pfet_05v0 L=6e-07 W=1.134e-05 AD=2.9484e-12 AS=4.9896e-12 PD=1.238e-05 PS=2.444e-05 NRD=0.0917108 NRS=0.155203 m=1 nf=2 $X=242235 $Y=57810 $D=8
M894 281 808 VDD VDD pfet_05v0 L=1e-06 W=9e-07 AD=3.96e-13 AS=3.96e-13 PD=2.68e-06 PS=2.68e-06 NRD=0.488889 NRS=0.488889 m=1 nf=1 $X=243265 $Y=42525 $D=8
M895 CEN 617 619 VDD pfet_05v0 L=6e-07 W=2.27e-06 AD=9.988e-13 AS=9.988e-13 PD=5.42e-06 PS=5.42e-06 NRD=0.193833 NRS=0.193833 m=1 nf=1 $X=245925 $Y=59010 $D=8
M896 618 802 619 VDD pfet_05v0 L=6e-07 W=9.6e-07 AD=4.224e-13 AS=4.224e-13 PD=2.8e-06 PS=2.8e-06 NRD=0.458333 NRS=0.458333 m=1 nf=1 $X=245925 $Y=64875 $D=8
M897 317 281 VDD VDD pfet_05v0 L=6e-07 W=1.89e-06 AD=8.316e-13 AS=8.316e-13 PD=4.66e-06 PS=4.66e-06 NRD=0.232804 NRS=0.232804 m=1 nf=1 $X=246495 $Y=41535 $D=8
M898 354 317 VDD VDD pfet_05v0 L=6e-07 W=7.54e-06 AD=1.9604e-12 AS=3.3176e-12 PD=8.58e-06 PS=1.684e-05 NRD=0.137931 NRS=0.233422 m=1 nf=2 $X=249065 $Y=39655 $D=8
M899 250 468 VDD VDD pfet_05v0 L=6e-07 W=0.0001248 AD=3.2448e-11 AS=3.69283e-11 PD=0.00013 PS=0.000130718 NRD=0.208333 NRS=0.237099 m=1 nf=10 $X=240535 $Y=94430 $D=8
M900 445 354 VDD VDD pfet_05v0 L=6e-07 W=1.95e-05 AD=5.07e-12 AS=8.58e-12 PD=2.002e-05 PS=3.988e-05 NRD=0.0133333 NRS=0.0225641 m=1 nf=1 $X=256125 $Y=53590 $D=8
M901 VDD CLK 445 VDD pfet_05v0 L=6e-07 W=1.95e-05 AD=0 AS=0 PD=0 PS=0 NRD=0 NRS=0 m=1 nf=1 $X=257245 $Y=53590 $D=8
M902 445 616 VDD VDD pfet_05v0 L=6e-07 W=1.95e-05 AD=8.58e-12 AS=5.07e-12 PD=3.988e-05 PS=2.002e-05 NRD=0.0225641 NRS=0.0133333 m=1 nf=1 $X=258365 $Y=53590 $D=8
M903 VDD 495 468 VDD pfet_05v0 L=6e-07 W=2.268e-05 AD=5.8968e-12 AS=9.9792e-12 PD=2.32e-05 PS=4.624e-05 NRD=0.0114638 NRS=0.0194004 m=1 nf=1 $X=262120 $Y=50420 $D=8
M904 468 445 VDD VDD pfet_05v0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.64e-05 PS=4.64e-05 NRD=0.0229277 NRS=0.0229277 m=1 nf=2 $X=263240 $Y=50420 $D=8
M905 468 495 VDD VDD pfet_05v0 L=6e-07 W=2.268e-05 AD=9.9792e-12 AS=5.8968e-12 PD=4.624e-05 PS=2.32e-05 NRD=0.0194004 NRS=0.0114638 m=1 nf=1 $X=265480 $Y=50420 $D=8
M906 VDD 468 495 VDD pfet_05v0 L=6e-07 W=2.268e-05 AD=5.8968e-12 AS=9.9792e-12 PD=2.32e-05 PS=4.624e-05 NRD=0.0114638 NRS=0.0194004 m=1 nf=1 $X=268545 $Y=50420 $D=8
M907 495 607 VDD VDD pfet_05v0 L=6e-07 W=4.536e-05 AD=1.17936e-11 AS=1.17936e-11 PD=4.64e-05 PS=4.64e-05 NRD=0.0229277 NRS=0.0229277 m=1 nf=2 $X=269665 $Y=50420 $D=8
M908 495 468 VDD VDD pfet_05v0 L=6e-07 W=2.268e-05 AD=9.9792e-12 AS=5.8968e-12 PD=4.624e-05 PS=2.32e-05 NRD=0.0194004 NRS=0.0114638 m=1 nf=1 $X=271905 $Y=50420 $D=8
M909 1 250 VDD VDD pfet_05v0 L=6e-07 W=0.0003674 AD=9.5524e-11 AS=1.02119e-10 PD=0.0003778 PS=0.000378518 NRD=0.28307 NRS=0.302613 m=1 nf=20 $X=253180 $Y=88540 $D=8
M910 VDD VSS VDD VDD pfet_05v0 L=3.94e-06 W=0.000181335 AD=0 AS=1.05339e-10 PD=0 PS=0.000412 NRD=0 NRS=3.48863 m=1 nf=33 $X=273750 $Y=180915 $D=8
M911 VDD 4304 4305 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=179690 $D=8
M912 VDD 5383 5384 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=180970 $D=8
M913 VDD 5385 5386 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=197690 $D=8
M914 VDD 5387 5388 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=198970 $D=8
M915 VDD 5389 5390 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=215690 $D=8
M916 VDD 5391 5392 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=216970 $D=8
M917 VDD 5393 5394 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=233690 $D=8
M918 VDD 5395 5396 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=234970 $D=8
M919 VDD 5397 5398 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=251690 $D=8
M920 VDD 5399 5400 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=252970 $D=8
M921 VDD 5401 5402 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=269690 $D=8
M922 VDD 5403 5404 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=270970 $D=8
M923 VDD 5405 5406 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=287690 $D=8
M924 VDD 5407 5408 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=288970 $D=8
M925 VDD 5409 5410 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=305690 $D=8
M926 VDD 5411 5412 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=306970 $D=8
M927 VDD 5413 5414 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=323690 $D=8
M928 VDD 4306 4307 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=304720 $Y=324970 $D=8
M929 4304 4305 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=179690 $D=8
M930 5383 5384 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=180970 $D=8
M931 5385 5386 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=197690 $D=8
M932 5387 5388 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=198970 $D=8
M933 5389 5390 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=215690 $D=8
M934 5391 5392 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=216970 $D=8
M935 5393 5394 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=233690 $D=8
M936 5395 5396 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=234970 $D=8
M937 5397 5398 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=251690 $D=8
M938 5399 5400 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=252970 $D=8
M939 5401 5402 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=269690 $D=8
M940 5403 5404 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=270970 $D=8
M941 5405 5406 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=287690 $D=8
M942 5407 5408 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=288970 $D=8
M943 5409 5410 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=305690 $D=8
M944 5411 5412 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=306970 $D=8
M945 5413 5414 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=323690 $D=8
M946 4306 4307 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=305860 $Y=324970 $D=8
M947 VDD 4281 4283 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=179690 $D=8
M948 VDD 5416 5415 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=310720 $Y=180970 $D=8
M949 4281 4283 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=179690 $D=8
M950 5416 5415 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=311860 $Y=180970 $D=8
M951 4644 4099 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=311500 $Y=160970 $D=8
M952 4645 4099 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=311500 $Y=164845 $D=8
M953 4793 4573 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=311715 $Y=112830 $D=8
M954 VDD 4277 4279 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=179690 $D=8
M955 VDD 5418 5417 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=313720 $Y=180970 $D=8
M956 4277 4279 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=179690 $D=8
M957 5418 5417 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=314860 $Y=180970 $D=8
M958 4794 4574 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=314245 $Y=112830 $D=8
M959 4647 4099 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=314600 $Y=160970 $D=8
M960 4646 4099 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=314600 $Y=164845 $D=8
M961 VDD 4273 4275 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=179690 $D=8
M962 VDD 5420 5419 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=316720 $Y=180970 $D=8
M963 4273 4275 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=179690 $D=8
M964 5420 5419 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=317860 $Y=180970 $D=8
M965 4648 4099 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=317695 $Y=160970 $D=8
M966 4649 4099 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=317695 $Y=164845 $D=8
M967 4795 4575 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=317910 $Y=112830 $D=8
M968 VDD 4269 4271 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=179690 $D=8
M969 VDD 5422 5421 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=319720 $Y=180970 $D=8
M970 4269 4271 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=179690 $D=8
M971 5422 5421 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=320860 $Y=180970 $D=8
M972 4796 4576 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=320440 $Y=112830 $D=8
M973 4651 4099 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=320795 $Y=160970 $D=8
M974 4650 4099 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=320795 $Y=164845 $D=8
M975 VDD 4209 4211 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=179690 $D=8
M976 VDD 5424 5423 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=322720 $Y=180970 $D=8
M977 4209 4211 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=179690 $D=8
M978 5424 5423 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=323860 $Y=180970 $D=8
M979 4652 4099 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=323885 $Y=160970 $D=8
M980 4653 4099 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=323885 $Y=164845 $D=8
M981 4797 4577 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=324100 $Y=112830 $D=8
M982 VDD 4205 4207 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=179690 $D=8
M983 VDD 5426 5425 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=325720 $Y=180970 $D=8
M984 4205 4207 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=179690 $D=8
M985 5426 5425 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=326860 $Y=180970 $D=8
M986 4798 4578 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=326630 $Y=112830 $D=8
M987 4655 4099 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=326985 $Y=160970 $D=8
M988 4654 4099 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=326985 $Y=164845 $D=8
M989 VDD 4217 4219 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=179690 $D=8
M990 VDD 5428 5427 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=328720 $Y=180970 $D=8
M991 4217 4219 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=179690 $D=8
M992 5428 5427 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=329860 $Y=180970 $D=8
M993 4656 4099 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=330080 $Y=160970 $D=8
M994 4657 4099 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=330080 $Y=164845 $D=8
M995 4799 4579 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=330295 $Y=112830 $D=8
M996 VDD 4213 4215 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=179690 $D=8
M997 VDD 5430 5429 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=331720 $Y=180970 $D=8
M998 4213 4215 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=179690 $D=8
M999 5430 5429 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=332860 $Y=180970 $D=8
M1000 4737 4580 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=332825 $Y=112830 $D=8
M1001 886 4099 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=333000 $Y=160970 $D=8
M1002 887 4099 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=333000 $Y=164845 $D=8
M1003 900 898 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=336455 $Y=160970 $D=8
M1004 901 898 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=336455 $Y=164845 $D=8
M1005 VDD 4529 4531 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=179690 $D=8
M1006 VDD 5449 5450 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=337720 $Y=180970 $D=8
M1007 4741 4573 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=336500 $Y=112830 $D=8
M1008 4529 4531 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=179690 $D=8
M1009 5449 5450 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=338860 $Y=180970 $D=8
M1010 5339 4574 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=339025 $Y=112830 $D=8
M1011 4712 898 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=339380 $Y=160970 $D=8
M1012 4713 898 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=339380 $Y=164845 $D=8
M1013 VDD 4525 4527 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=179690 $D=8
M1014 VDD 5447 5448 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=340720 $Y=180970 $D=8
M1015 4525 4527 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=179690 $D=8
M1016 5447 5448 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=341860 $Y=180970 $D=8
M1017 4711 898 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=342475 $Y=160970 $D=8
M1018 4710 898 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=342475 $Y=164845 $D=8
M1019 VDD 4521 4523 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=179690 $D=8
M1020 VDD 5453 5454 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=343720 $Y=180970 $D=8
M1021 5338 4575 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=342690 $Y=112830 $D=8
M1022 4521 4523 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=179690 $D=8
M1023 5453 5454 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=344860 $Y=180970 $D=8
M1024 5337 4576 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=345220 $Y=112830 $D=8
M1025 4708 898 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=345575 $Y=160970 $D=8
M1026 4709 898 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=345575 $Y=164845 $D=8
M1027 VDD 4517 4519 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=179690 $D=8
M1028 VDD 5451 5452 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=346720 $Y=180970 $D=8
M1029 4517 4519 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=179690 $D=8
M1030 5451 5452 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=347860 $Y=180970 $D=8
M1031 VDD 4513 4515 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=179690 $D=8
M1032 VDD 5457 5458 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=349720 $Y=180970 $D=8
M1033 4707 898 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=348665 $Y=160970 $D=8
M1034 4706 898 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=348665 $Y=164845 $D=8
M1035 5336 4577 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=348880 $Y=112830 $D=8
M1036 4513 4515 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=179690 $D=8
M1037 5457 5458 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=350860 $Y=180970 $D=8
M1038 5335 4578 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=351410 $Y=112830 $D=8
M1039 VDD 4509 4511 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=179690 $D=8
M1040 VDD 5455 5456 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=352720 $Y=180970 $D=8
M1041 4704 898 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=351765 $Y=160970 $D=8
M1042 4705 898 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=351765 $Y=164845 $D=8
M1043 4509 4511 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=179690 $D=8
M1044 5455 5456 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=353860 $Y=180970 $D=8
M1045 VDD 4505 4507 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=179690 $D=8
M1046 VDD 5461 5462 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=355720 $Y=180970 $D=8
M1047 4703 898 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=354860 $Y=160970 $D=8
M1048 4702 898 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=354860 $Y=164845 $D=8
M1049 5334 4579 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=355075 $Y=112830 $D=8
M1050 4505 4507 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=179690 $D=8
M1051 5461 5462 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=356860 $Y=180970 $D=8
M1052 VDD 4501 4503 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=179690 $D=8
M1053 VDD 5459 5460 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=358720 $Y=180970 $D=8
M1054 5333 4580 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=357605 $Y=112830 $D=8
M1055 4700 898 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=357960 $Y=160970 $D=8
M1056 4701 898 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=357960 $Y=164845 $D=8
M1057 4501 4503 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=179690 $D=8
M1058 5459 5460 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=359860 $Y=180970 $D=8
M1059 VDD 4297 4299 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=179690 $D=8
M1060 VDD 5432 5431 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=364720 $Y=180970 $D=8
M1061 4297 4299 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=179690 $D=8
M1062 5432 5431 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=365860 $Y=180970 $D=8
M1063 4658 4100 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=365500 $Y=160970 $D=8
M1064 4659 4100 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=365500 $Y=164845 $D=8
M1065 4800 4573 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=365715 $Y=112830 $D=8
M1066 VDD 4293 4295 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=179690 $D=8
M1067 VDD 5434 5433 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=367720 $Y=180970 $D=8
M1068 4293 4295 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=179690 $D=8
M1069 5434 5433 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=368860 $Y=180970 $D=8
M1070 4801 4574 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=368245 $Y=112830 $D=8
M1071 4661 4100 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=368600 $Y=160970 $D=8
M1072 4660 4100 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=368600 $Y=164845 $D=8
M1073 VDD 4289 4291 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=179690 $D=8
M1074 VDD 5436 5435 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=370720 $Y=180970 $D=8
M1075 4289 4291 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=179690 $D=8
M1076 5436 5435 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=371860 $Y=180970 $D=8
M1077 4662 4100 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=371695 $Y=160970 $D=8
M1078 4663 4100 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=371695 $Y=164845 $D=8
M1079 4802 4575 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=371910 $Y=112830 $D=8
M1080 VDD 4285 4287 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=179690 $D=8
M1081 VDD 5438 5437 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=373720 $Y=180970 $D=8
M1082 4285 4287 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=179690 $D=8
M1083 5438 5437 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=374860 $Y=180970 $D=8
M1084 4803 4576 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=374440 $Y=112830 $D=8
M1085 4665 4100 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=374795 $Y=160970 $D=8
M1086 4664 4100 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=374795 $Y=164845 $D=8
M1087 VDD 4225 4227 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=179690 $D=8
M1088 VDD 5440 5439 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=376720 $Y=180970 $D=8
M1089 4225 4227 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=179690 $D=8
M1090 5440 5439 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=377860 $Y=180970 $D=8
M1091 4666 4100 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=377885 $Y=160970 $D=8
M1092 4667 4100 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=377885 $Y=164845 $D=8
M1093 4804 4577 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=378100 $Y=112830 $D=8
M1094 VDD 4221 4223 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=179690 $D=8
M1095 VDD 5442 5441 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=379720 $Y=180970 $D=8
M1096 4221 4223 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=179690 $D=8
M1097 5442 5441 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=380860 $Y=180970 $D=8
M1098 4805 4578 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=380630 $Y=112830 $D=8
M1099 4669 4100 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=380985 $Y=160970 $D=8
M1100 4668 4100 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=380985 $Y=164845 $D=8
M1101 VDD 4233 4235 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=179690 $D=8
M1102 VDD 5444 5443 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=382720 $Y=180970 $D=8
M1103 4233 4235 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=179690 $D=8
M1104 5444 5443 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=383860 $Y=180970 $D=8
M1105 4670 4100 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=384080 $Y=160970 $D=8
M1106 4671 4100 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=384080 $Y=164845 $D=8
M1107 4806 4579 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=384295 $Y=112830 $D=8
M1108 VDD 4229 4231 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=179690 $D=8
M1109 VDD 5446 5445 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=385720 $Y=180970 $D=8
M1110 4229 4231 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=179690 $D=8
M1111 5446 5445 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=386860 $Y=180970 $D=8
M1112 4738 4580 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=386825 $Y=112830 $D=8
M1113 889 4100 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=387000 $Y=160970 $D=8
M1114 890 4100 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=387000 $Y=164845 $D=8
M1115 903 879 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=390455 $Y=160970 $D=8
M1116 904 879 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.79025e-12 AS=4.99565e-12 PD=7.87e-06 PS=9.75e-06 NRD=0.153959 NRS=0.429619 m=1 nf=2 $X=390455 $Y=164845 $D=8
M1117 VDD 4561 4563 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=179690 $D=8
M1118 VDD 5465 5466 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=391720 $Y=180970 $D=8
M1119 4742 4573 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.72675e-13 AS=1.84882e-12 PD=4.28e-06 PS=5.46e-06 NRD=0.441077 NRS=0.838384 m=1 nf=2 $X=390500 $Y=112830 $D=8
M1120 4561 4563 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=179690 $D=8
M1121 5465 5466 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=392860 $Y=180970 $D=8
M1122 5346 4574 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=393025 $Y=112830 $D=8
M1123 4726 879 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=393380 $Y=160970 $D=8
M1124 4727 879 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.39037e-12 PD=7.86e-06 PS=9.395e-06 NRD=0.152493 NRS=0.377566 m=1 nf=2 $X=393380 $Y=164845 $D=8
M1125 VDD 4557 4559 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=179690 $D=8
M1126 VDD 5463 5464 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=394720 $Y=180970 $D=8
M1127 4557 4559 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=179690 $D=8
M1128 5463 5464 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=395860 $Y=180970 $D=8
M1129 4725 879 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=396475 $Y=160970 $D=8
M1130 4724 879 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=396475 $Y=164845 $D=8
M1131 VDD 4553 4555 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=179690 $D=8
M1132 VDD 5469 5470 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=397720 $Y=180970 $D=8
M1133 5345 4575 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=396690 $Y=112830 $D=8
M1134 4553 4555 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=179690 $D=8
M1135 5469 5470 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=398860 $Y=180970 $D=8
M1136 5344 4576 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=399220 $Y=112830 $D=8
M1137 4722 879 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=399575 $Y=160970 $D=8
M1138 4723 879 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=399575 $Y=164845 $D=8
M1139 VDD 4549 4551 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=179690 $D=8
M1140 VDD 5467 5468 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=400720 $Y=180970 $D=8
M1141 4549 4551 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=179690 $D=8
M1142 5467 5468 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=401860 $Y=180970 $D=8
M1143 VDD 4545 4547 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=179690 $D=8
M1144 VDD 5473 5474 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=403720 $Y=180970 $D=8
M1145 4721 879 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=402665 $Y=160970 $D=8
M1146 4720 879 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.68875e-12 PD=7.86e-06 PS=9.57e-06 NRD=0.152493 NRS=0.403226 m=1 nf=2 $X=402665 $Y=164845 $D=8
M1147 5343 4577 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83397e-12 PD=4.29e-06 PS=5.44e-06 NRD=0.444444 NRS=0.83165 m=1 nf=2 $X=402880 $Y=112830 $D=8
M1148 4545 4547 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=179690 $D=8
M1149 5473 5474 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=404860 $Y=180970 $D=8
M1150 5342 4578 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=405410 $Y=112830 $D=8
M1151 VDD 4541 4543 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=179690 $D=8
M1152 VDD 5471 5472 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=406720 $Y=180970 $D=8
M1153 4718 879 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=405765 $Y=160970 $D=8
M1154 4719 879 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=405765 $Y=164845 $D=8
M1155 4541 4543 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=179690 $D=8
M1156 5471 5472 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=407860 $Y=180970 $D=8
M1157 VDD 4537 4539 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=179690 $D=8
M1158 VDD 5477 5478 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=409720 $Y=180970 $D=8
M1159 4717 879 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=408860 $Y=160970 $D=8
M1160 4716 879 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=4.69727e-12 PD=7.86e-06 PS=9.575e-06 NRD=0.152493 NRS=0.403959 m=1 nf=2 $X=408860 $Y=164845 $D=8
M1161 5341 4579 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.83769e-12 PD=4.29e-06 PS=5.445e-06 NRD=0.444444 NRS=0.833333 m=1 nf=2 $X=409075 $Y=112830 $D=8
M1162 4537 4539 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=179690 $D=8
M1163 5477 5478 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=410860 $Y=180970 $D=8
M1164 VDD 4533 4535 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=179690 $D=8
M1165 VDD 5475 5476 VDD pfet_05v0 L=6e-07 W=6e-07 AD=8.52e-13 AS=2.7e-13 PD=5.32e-06 PS=2.1e-06 NRD=2.36667 NRS=0.75 m=1 nf=1 $X=412720 $Y=180970 $D=8
M1166 5340 4580 VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=1.8414e-12 PD=4.29e-06 PS=6.935e-06 NRD=0.444444 NRS=0.835017 m=1 nf=2 $X=411605 $Y=112830 $D=8
M1167 4714 879 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=411960 $Y=160970 $D=8
M1168 4715 879 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=5.2173e-12 PD=7.86e-06 PS=1.329e-05 NRD=0.152493 NRS=0.44868 m=1 nf=2 $X=411960 $Y=164845 $D=8
M1169 VDD VSS VDD VDD pfet_05v0 L=2.365e-06 W=8.19e-05 AD=0 AS=6.1309e-11 PD=0 PS=0.000217698 NRD=0 NRS=11.8457 m=1 nf=36 $X=303025 $Y=171065 $D=8
M1170 4533 4535 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=179690 $D=8
M1171 5475 5476 VDD VDD pfet_05v0 L=6e-07 W=6e-07 AD=2.7e-13 AS=8.52e-13 PD=2.1e-06 PS=5.32e-06 NRD=0.75 NRS=2.36667 m=1 nf=1 $X=413860 $Y=180970 $D=8
M1172 614 879 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=6.35965e-12 PD=7.86e-06 PS=1.737e-05 NRD=0.152493 NRS=0.546921 m=1 nf=2 $X=418655 $Y=160970 $D=8
M1173 615 879 VDD VDD pfet_05v0 L=6e-07 W=6.82e-06 AD=1.7732e-12 AS=6.35965e-12 PD=7.86e-06 PS=1.737e-05 NRD=0.152493 NRS=0.546921 m=1 nf=2 $X=418655 $Y=164845 $D=8
M1174 606 614 VDD VDD pfet_05v0 L=6e-07 W=7.02e-06 AD=1.8252e-12 AS=3.0888e-12 PD=8.06e-06 PS=1.58e-05 NRD=0.148148 NRS=0.250712 m=1 nf=2 $X=418770 $Y=97440 $D=8
M1175 607 606 VDD VDD pfet_05v0 L=6e-07 W=2.128e-05 AD=5.5328e-12 AS=9.3632e-12 PD=2.232e-05 PS=4.432e-05 NRD=0.0488722 NRS=0.0827068 m=1 nf=2 $X=418790 $Y=67070 $D=8
M1176 613 VDD VDD VDD pfet_05v0 L=6e-07 W=2.97e-06 AD=9.801e-13 AS=2.33887e-12 PD=4.29e-06 PS=9.09e-06 NRD=0.444444 NRS=1.06061 m=1 nf=2 $X=418870 $Y=112830 $D=8
X1185 614 614 613 VDD pfet_05v0_I09 $T=419815 124190 0 180 $X=418175 $Y=116760
X1186 615 615 613 VDD pfet_05v0_I09 $T=419815 151940 0 180 $X=418175 $Y=144510
X1187 615 614 879 VDD pfet_05v0_I09 $T=419825 159875 0 180 $X=418185 $Y=152445
X1188 614 614 VDD VSS nfet_05v0_I12 $T=419815 133465 0 180 $X=418535 $Y=126035
X1189 615 615 VDD VSS nfet_05v0_I12 $T=419815 143485 0 180 $X=418535 $Y=136055
X1195 VDD 618 616 pmos_1p2$$46273580 $T=242390 65835 1 0 $X=240960 $Y=64015
X1196 VSS 617 802 VSS nmos_1p2$$46563372 $T=233925 66830 0 0 $X=232780 $Y=66145
X1197 618 VSS 616 VSS nmos_1p2$$46563372 $T=243510 68190 1 0 $X=242365 $Y=66555
X1198 619 618 617 VSS nmos_1p2$$46563372 $T=246080 68190 1 0 $X=244935 $Y=66555
X1200 880 VSS Q[0] D[0] 4097 1 VDD 881 882 WEN[0] 4616 4617 4618 4619 4620 4621 4622 4623 4624 4625
+ 4626 4627 4628 4629 4735 870 4571 4570 4569 4568 4567 4566 4565 4564 4572 4779 4780 4781 4782 4783
+ 4784 4785
+ saout_m2 $T=9775 25090 0 0 $X=8430 $Y=7315
X1201 864 VSS Q[2] D[2] 4098 1 VDD 883 884 WEN[2] 4630 4631 4632 4633 4634 4635 4636 4637 4638 4639
+ 4640 4641 4642 4643 4736 870 4571 4570 4569 4568 4567 4566 4565 4564 4572 4786 4787 4788 4789 4790
+ 4791 4792
+ saout_m2 $T=63775 25090 0 0 $X=62430 $Y=7315
X1202 885 VSS Q[4] D[4] 4099 1 VDD 886 887 WEN[4] 4644 4645 4646 4647 4648 4649 4650 4651 4652 4653
+ 4654 4655 4656 4657 4737 870 4573 4574 4575 4576 4577 4578 4579 4580 4572 4793 4794 4795 4796 4797
+ 4798 4799
+ saout_m2 $T=307655 25090 0 0 $X=306310 $Y=7315
X1203 888 VSS Q[6] D[6] 4100 1 VDD 889 890 WEN[6] 4658 4659 4660 4661 4662 4663 4664 4665 4666 4667
+ 4668 4669 4670 4671 4738 870 4573 4574 4575 4576 4577 4578 4579 4580 4572 4800 4801 4802 4803 4804
+ 4805 4806
+ saout_m2 $T=361655 25090 0 0 $X=360310 $Y=7315
X1204 VSS VSS 4172 4173 4174 4175 4176 4177 4178 4179 ICV_6 $T=27210 176130 1 180 $X=23870 $Y=175790
X1205 VSS VSS 4180 4181 4182 4183 4184 4185 4186 4187 ICV_6 $T=33210 176130 1 180 $X=29870 $Y=175790
X1206 VSS VSS 4188 4189 4190 4191 4192 4193 4194 4195 ICV_6 $T=81210 176130 1 180 $X=77870 $Y=175790
X1207 VSS VSS 4196 4197 4198 4199 4200 4201 4202 4203 ICV_6 $T=87210 176130 1 180 $X=83870 $Y=175790
X1208 VSS VSS 4204 4205 4206 4207 4208 4209 4210 4211 ICV_6 $T=325090 176130 1 180 $X=321750 $Y=175790
X1209 VSS VSS 4212 4213 4214 4215 4216 4217 4218 4219 ICV_6 $T=331090 176130 1 180 $X=327750 $Y=175790
X1210 VSS VSS 4220 4221 4222 4223 4224 4225 4226 4227 ICV_6 $T=379090 176130 1 180 $X=375750 $Y=175790
X1211 VSS VSS 4228 4229 4230 4231 4232 4233 4234 4235 ICV_6 $T=385090 176130 1 180 $X=381750 $Y=175790
X1218 VSS 4236 4237 4238 4239 4240 4241 4242 4243 4244 4245 4246 4247 4248 4249 4250 4251 ICV_14 $T=12210 176130 1 180 $X=8870 $Y=175790
X1219 VSS 4252 4253 4254 4255 4256 4257 4258 4259 4260 4261 4262 4263 4264 4265 4266 4267 ICV_14 $T=66210 176130 1 180 $X=62870 $Y=175790
X1220 VSS 4268 4269 4270 4271 4272 4273 4274 4275 4276 4277 4278 4279 4280 4281 4282 4283 ICV_14 $T=310090 176130 1 180 $X=306750 $Y=175790
X1221 VSS 4284 4285 4286 4287 4288 4289 4290 4291 4292 4293 4294 4295 4296 4297 4298 4299 ICV_14 $T=364090 176130 1 180 $X=360750 $Y=175790
X1226 VDD VSS 4101 4102 4103 4104 4105 4106 4107 4108 4672 4673 4674 4675 4676 4677 4678 4679 4680 4681
+ 4682 4683 4684 4685 894 893 4624 4625 4626 4627 4628 4629 882 881 4616 4617 4618 4619 4620 4621
+ 4622 4623 4807 4808 4809 4810 4811 4812 4813 4814 4815 4816 4817 4818 4819 4820 4821 4822 4823 4824
+ 4825 4826 4827 4828 4829 4830 4831 4832 4833 4834 4835 4836 4837 4838 4839 4840 4841 4842 4843 4844
+ 4845 4846 4847 4848 4849 4850 4851 4852 4853 4854 4855 4856 4857 4858 4859 4860 4861 4862 4863 4864
+ 4865 4866 4867 4868 4869 4870
+ ICV_35 $T=12210 185130 1 180 $X=8870 $Y=180290
X1227 VDD VSS 4109 4110 4111 4112 4113 4114 4115 4116 4672 4673 4674 4675 4676 4677 4678 4679 4680 4681
+ 4682 4683 4684 4685 894 893 4624 4625 4626 4627 4628 4629 882 881 4616 4617 4618 4619 4620 4621
+ 4622 4623 4871 4872 4873 4874 4875 4876 4877 4878 4879 4880 4881 4882 4883 4884 4885 4886 4887 4888
+ 4889 4890 4891 4892 4893 4894 4895 4896 4897 4898 4899 4900 4901 4902 4903 4904 4905 4906 4907 4908
+ 4909 4910 4911 4912 4913 4914 4915 4916 4917 4918 4919 4920 4921 4922 4923 4924 4925 4926 4927 4928
+ 4929 4930 4931 4932 4933 4934
+ ICV_35 $T=12210 221130 1 180 $X=8870 $Y=216290
X1228 VDD VSS 4117 4118 4119 4120 4121 4122 4123 4124 4672 4673 4674 4675 4676 4677 4678 4679 4680 4681
+ 4682 4683 4684 4685 894 893 4624 4625 4626 4627 4628 4629 882 881 4616 4617 4618 4619 4620 4621
+ 4622 4623 4935 4936 4937 4938 4939 4940 4941 4942 4943 4944 4945 4946 4947 4948 4949 4950 4951 4952
+ 4953 4954 4955 4956 4957 4958 4959 4960 4961 4962 4963 4964 4965 4966 4967 4968 4969 4970 4971 4972
+ 4973 4974 4975 4976 4977 4978 4979 4980 4981 4982 4983 4984 4985 4986 4987 4988 4989 4990 4991 4992
+ 4993 4994 4995 4996 4997 4998
+ ICV_35 $T=12210 257130 1 180 $X=8870 $Y=252290
X1229 VDD VSS 4125 4126 4127 4128 4129 4130 4131 4132 4672 4673 4674 4675 4676 4677 4678 4679 4680 4681
+ 4682 4683 4684 4685 894 893 4624 4625 4626 4627 4628 4629 882 881 4616 4617 4618 4619 4620 4621
+ 4622 4623 4999 5000 5001 5002 5003 5004 5005 5006 5007 5008 5009 5010 5011 5012 5013 5014 5015 5016
+ 5017 5018 5019 5020 5021 5022 5023 5024 5025 5026 5027 5028 5029 5030 5031 5032 5033 5034 5035 5036
+ 5037 5038 5039 5040 5041 5042 5043 5044 5045 5046 5047 5048 5049 5050 5051 5052 5053 5054 5055 5056
+ 5057 5058 5059 5060 5061 5062
+ ICV_35 $T=12210 293130 1 180 $X=8870 $Y=288290
X1230 VDD VSS 4101 4102 4103 4104 4105 4106 4107 4108 4686 4687 4688 4689 4690 4691 4692 4693 4694 4695
+ 4696 4697 4698 4699 897 896 4638 4639 4640 4641 4642 4643 884 883 4630 4631 4632 4633 4634 4635
+ 4636 4637 5063 5064 5065 5066 5067 5068 5069 5070 5071 5072 5073 5074 5075 5076 5077 5078 5079 5080
+ 5081 5082 5083 5084 5085 5086 5087 5088 5089 5090 5091 5092 5093 5094 5095 5096 5097 5098 5099 5100
+ 5101 5102 5103 5104 5105 5106 5107 5108 5109 5110 5111 5112 5113 5114 5115 5116 5117 5118 5119 5120
+ 5121 5122 5123 5124 5125 5126
+ ICV_35 $T=66210 185130 1 180 $X=62870 $Y=180290
X1231 VDD VSS 4109 4110 4111 4112 4113 4114 4115 4116 4686 4687 4688 4689 4690 4691 4692 4693 4694 4695
+ 4696 4697 4698 4699 897 896 4638 4639 4640 4641 4642 4643 884 883 4630 4631 4632 4633 4634 4635
+ 4636 4637 5127 5128 5129 5130 5131 5132 5133 5134 5135 5136 5137 5138 5139 5140 5141 5142 5143 5144
+ 5145 5146 5147 5148 5149 5150 5151 5152 5153 5154 5155 5156 5157 5158 5159 5160 5161 5162 5163 5164
+ 5165 5166 5167 5168 5169 5170 5171 5172 5173 5174 5175 5176 5177 5178 5179 5180 5181 5182 5183 5184
+ 5185 5186 5187 5188 5189 5190
+ ICV_35 $T=66210 221130 1 180 $X=62870 $Y=216290
X1232 VDD VSS 4117 4118 4119 4120 4121 4122 4123 4124 4686 4687 4688 4689 4690 4691 4692 4693 4694 4695
+ 4696 4697 4698 4699 897 896 4638 4639 4640 4641 4642 4643 884 883 4630 4631 4632 4633 4634 4635
+ 4636 4637 5191 5192 5193 5194 5195 5196 5197 5198 5199 5200 5201 5202 5203 5204 5205 5206 5207 5208
+ 5209 5210 5211 5212 5213 5214 5215 5216 5217 5218 5219 5220 5221 5222 5223 5224 5225 5226 5227 5228
+ 5229 5230 5231 5232 5233 5234 5235 5236 5237 5238 5239 5240 5241 5242 5243 5244 5245 5246 5247 5248
+ 5249 5250 5251 5252 5253 5254
+ ICV_35 $T=66210 257130 1 180 $X=62870 $Y=252290
X1233 VDD VSS 4125 4126 4127 4128 4129 4130 4131 4132 4686 4687 4688 4689 4690 4691 4692 4693 4694 4695
+ 4696 4697 4698 4699 897 896 4638 4639 4640 4641 4642 4643 884 883 4630 4631 4632 4633 4634 4635
+ 4636 4637 5255 5256 5257 5258 5259 5260 5261 5262 5263 5264 5265 5266 5267 5268 5269 5270 5271 5272
+ 5273 5274 5275 5276 5277 5278 5279 5280 5281 5282 5283 5284 5285 5286 5287 5288 5289 5290 5291 5292
+ 5293 5294 5295 5296 5297 5298 5299 5300 5301 5302 5303 5304 5305 5306 5307 5308 5309 5310 5311 5312
+ 5313 5314 5315 5316 5317 5318
+ ICV_35 $T=66210 293130 1 180 $X=62870 $Y=288290
X1234 VSS 4308 4309 4310 4311 4312 4313 4314 4315 4316 4317 4318 4319 4320 4321 4322 4323 4324 4325 4326
+ 4327 4328 4329 4330 4331 4332 4333 4334 4335 4336 4337 4338 4339
+ ICV_15 $T=12210 329130 0 180 $X=8870 $Y=324290
X1235 VSS 4340 4341 4342 4343 4344 4345 4346 4347 4348 4349 4350 4351 4352 4353 4354 4355 4356 4357 4358
+ 4359 4360 4361 4362 4363 4364 4365 4366 4367 4368 4369 4370 4371
+ ICV_15 $T=39210 176130 1 180 $X=35870 $Y=175790
X1236 VSS 4372 4373 4374 4375 4376 4377 4378 4379 4380 4381 4382 4383 4384 4385 4386 4387 4388 4389 4390
+ 4391 4392 4393 4394 4395 4396 4397 4398 4399 4400 4401 4402 4403
+ ICV_15 $T=39210 329130 0 180 $X=35870 $Y=324290
X1237 VSS 4404 4405 4406 4407 4408 4409 4410 4411 4412 4413 4414 4415 4416 4417 4418 4419 4420 4421 4422
+ 4423 4424 4425 4426 4427 4428 4429 4430 4431 4432 4433 4434 4435
+ ICV_15 $T=66210 329130 0 180 $X=62870 $Y=324290
X1238 VSS 4436 4437 4438 4439 4440 4441 4442 4443 4444 4445 4446 4447 4448 4449 4450 4451 4452 4453 4454
+ 4455 4456 4457 4458 4459 4460 4461 4462 4463 4464 4465 4466 4467
+ ICV_15 $T=93210 176130 1 180 $X=89870 $Y=175790
X1239 VSS 4468 4469 4470 4471 4472 4473 4474 4475 4476 4477 4478 4479 4480 4481 4482 4483 4484 4485 4486
+ 4487 4488 4489 4490 4491 4492 4493 4494 4495 4496 4497 4498 4499
+ ICV_15 $T=93210 329130 0 180 $X=89870 $Y=324290
X1240 VSS 4500 4501 4502 4503 4504 4505 4506 4507 4508 4509 4510 4511 4512 4513 4514 4515 4516 4517 4518
+ 4519 4520 4521 4522 4523 4524 4525 4526 4527 4528 4529 4530 4531
+ ICV_15 $T=337090 176130 1 180 $X=333750 $Y=175790
X1241 VSS 4532 4533 4534 4535 4536 4537 4538 4539 4540 4541 4542 4543 4544 4545 4546 4547 4548 4549 4550
+ 4551 4552 4553 4554 4555 4556 4557 4558 4559 4560 4561 4562 4563
+ ICV_15 $T=391090 176130 1 180 $X=387750 $Y=175790
X1265 892 VSS Q[1] 891 D[1] 1 VDD 893 894 WEN[1] 4672 4673 4674 4675 4676 4677 4678 4679 4680 4681
+ 4682 4683 4684 4685 4739 870 4564 4565 4566 4567 4568 4569 4570 4571 4572 5319 5320 5321 5322 5323
+ 5324 5325
+ saout_R_m2 $T=65645 25125 1 180 $X=27480 $Y=6815
X1266 865 VSS Q[3] 895 D[3] 1 VDD 896 897 WEN[3] 4686 4687 4688 4689 4690 4691 4692 4693 4694 4695
+ 4696 4697 4698 4699 4740 870 4564 4565 4566 4567 4568 4569 4570 4571 4572 5326 5327 5328 5329 5330
+ 5331 5332
+ saout_R_m2 $T=119645 25125 1 180 $X=81480 $Y=6815
X1267 899 VSS Q[5] 898 D[5] 1 VDD 900 901 WEN[5] 4700 4701 4702 4703 4704 4705 4706 4707 4708 4709
+ 4710 4711 4712 4713 4741 870 4580 4579 4578 4577 4576 4575 4574 4573 4572 5333 5334 5335 5336 5337
+ 5338 5339
+ saout_R_m2 $T=363525 25125 1 180 $X=325360 $Y=6815
X1268 902 VSS Q[7] 879 D[7] 1 VDD 903 904 WEN[7] 4714 4715 4716 4717 4718 4719 4720 4721 4722 4723
+ 4724 4725 4726 4727 4742 870 4580 4579 4578 4577 4576 4575 4574 4573 4572 5340 5341 5342 5343 5344
+ 5345 5346
+ saout_R_m2 $T=417525 25125 1 180 $X=379360 $Y=6815
X1279 711 712 VSS 5347 5348 5349 5350 ICV_24 $T=123210 185130 0 180 $X=119870 $Y=180290
X1280 711 712 VSS 5351 5352 5353 5354 ICV_24 $T=123210 320130 0 180 $X=119870 $Y=315290
X1281 VDD VSS 711 712 5355 5356 5357 5358 ICV_25 $T=123210 194130 0 180 $X=119870 $Y=189290
X1282 VDD VSS 711 712 5359 5360 5361 5362 ICV_25 $T=123210 212130 0 180 $X=119870 $Y=207290
X1283 VDD VSS 711 712 5363 5364 5365 5366 ICV_25 $T=123210 230130 0 180 $X=119870 $Y=225290
X1284 VDD VSS 711 712 5367 5368 5369 5370 ICV_25 $T=123210 248130 0 180 $X=119870 $Y=243290
X1285 VDD VSS 711 712 5371 5372 5373 5374 ICV_25 $T=123210 266130 0 180 $X=119870 $Y=261290
X1286 VDD VSS 711 712 5375 5376 5377 5378 ICV_25 $T=123210 284130 0 180 $X=119870 $Y=279290
X1287 VDD VSS 711 712 5379 5380 5381 5382 ICV_25 $T=123210 302130 0 180 $X=119870 $Y=297290
X1305 VSS VDD 1 CLK VSS VSS 4589 4590 4594 4595 xpredec0 $T=146075 111460 0 0 $X=144630 $Y=111455
X1306 VSS VDD 1 CLK A[7] A[6] 4596 4597 4598 4599 xpredec0 $T=182970 111460 0 0 $X=181525 $Y=111455
X1311 VSS VDD 1 CLK 4570 4571 4564 4565 4566 4567 4568 4569 4580 4579 4578 4577 4576 4575 4574 4573
+ A[2] A[1] A[0]
+ ypredec1 $T=145470 26355 0 0 $X=146365 $Y=26735
X1312 VSS VDD 4596 4597 4598 4599 4600 4601 4602 4603 4604 4605 4606 4607 VDD 4101 4102 4103 4104 4105
+ 4106 4107 4108 4109 4110 4111 4112 4113 4114 4115 4116 4117 4118 4119 4120 4121 4122 4123 4124 4125
+ 4126 4127 4128 4129 4130 4131 4132 4134 4135 4136 4137 4138 4139 4140 4141 4142 4143 4144 4145 4146
+ 4147 4148 4149 4150 4151 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161 4162 4163 4164 4133 1
+ xdec32 $T=152015 180635 0 0 $X=152015 $Y=179495
X1315 803 VSS 805 nfet_05v0_I18 $T=175115 326995 0 90 $X=164385 $Y=326315
X1316 804 VSS 806 nfet_05v0_I18 $T=260115 326995 0 90 $X=249385 $Y=326315
X1320 VDD 803 805 pmos_1p2$$204216364 $T=189610 327150 0 90 $X=176320 $Y=325670
X1321 VDD 804 806 pmos_1p2$$204216364 $T=248135 327150 0 90 $X=234845 $Y=325670
X1322 805 VDD 2 VDD pfet_05v0_I01 $T=198405 326995 0 90 $X=191195 $Y=325955
X1323 1 2 VSS VDD pfet_05v0_I01 $T=219905 326995 0 90 $X=212695 $Y=325955
X1324 806 VDD 2 VDD pfet_05v0_I01 $T=233255 326995 0 90 $X=226045 $Y=325955
X1325 805 VSS 2 nfet_05v0_I04 $T=202950 326995 0 90 $X=199690 $Y=326315
X1326 806 VSS 2 nfet_05v0_I04 $T=224800 326995 0 90 $X=221540 $Y=326315
X1327 VSS VDD GWEN CLK 4572 870 wen_v2 $T=208415 16605 0 0 $X=208280 $Y=15275
X1328 VSS 1 VDD CLK A[5] A[4] A[3] 4600 4601 4602 4603 4604 4605 4606 4607 xpredec1 $T=219860 111460 0 0 $X=219855 $Y=111455
X1329 VDD 807 CLK pfet_05v0_I15 $T=234280 43425 1 0 $X=233240 $Y=41905
X1330 VDD 808 807 pfet_05v0_I15 $T=239670 43425 1 0 $X=238630 $Y=41905
X1331 VSS 807 CLK nfet_05v0_I16 $T=234280 46585 1 0 $X=233600 $Y=45365
X1332 VSS 808 807 nfet_05v0_I16 $T=239670 46585 1 0 $X=238990 $Y=45365
X1344 VDD VSS 713 714 5383 5384 5385 5386 ICV_18 $T=307090 180630 1 180 $X=303750 $Y=180290
X1345 VDD VSS 713 714 5387 5388 5389 5390 ICV_18 $T=307090 198630 1 180 $X=303750 $Y=198290
X1346 VDD VSS 713 714 5391 5392 5393 5394 ICV_18 $T=307090 216630 1 180 $X=303750 $Y=216290
X1347 VDD VSS 713 714 5395 5396 5397 5398 ICV_18 $T=307090 234630 1 180 $X=303750 $Y=234290
X1348 VDD VSS 713 714 5399 5400 5401 5402 ICV_18 $T=307090 252630 1 180 $X=303750 $Y=252290
X1349 VDD VSS 713 714 5403 5404 5405 5406 ICV_18 $T=307090 270630 1 180 $X=303750 $Y=270290
X1350 VDD VSS 713 714 5407 5408 5409 5410 ICV_18 $T=307090 288630 1 180 $X=303750 $Y=288290
X1351 VDD VSS 713 714 5411 5412 5413 5414 ICV_18 $T=307090 306630 1 180 $X=303750 $Y=306290
X1352 VSS VDD 804 4133 4134 4135 4136 4137 4138 4139 4140 4141 4142 4143 4144 4145 4146 4147 4148 4149
+ 4150 4151 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161 4162 4163 4164 4644 4645 4646 4647 5415
+ 5416 5417 5418
+ ICV_16 $T=310090 180630 0 0 $X=309750 $Y=180290
X1353 VSS VDD 804 4133 4134 4135 4136 4137 4138 4139 4140 4141 4142 4143 4144 4145 4146 4147 4148 4149
+ 4150 4151 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161 4162 4163 4164 4648 4649 4650 4651 5419
+ 5420 5421 5422
+ ICV_16 $T=316090 180630 0 0 $X=315750 $Y=180290
X1354 VSS VDD 804 4133 4134 4135 4136 4137 4138 4139 4140 4141 4142 4143 4144 4145 4146 4147 4148 4149
+ 4150 4151 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161 4162 4163 4164 4652 4653 4654 4655 5423
+ 5424 5425 5426
+ ICV_16 $T=322090 180630 0 0 $X=321750 $Y=180290
X1355 VSS VDD 804 4133 4134 4135 4136 4137 4138 4139 4140 4141 4142 4143 4144 4145 4146 4147 4148 4149
+ 4150 4151 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161 4162 4163 4164 4656 4657 887 886 5427
+ 5428 5429 5430
+ ICV_16 $T=328090 180630 0 0 $X=327750 $Y=180290
X1356 VSS VDD 804 4133 4134 4135 4136 4137 4138 4139 4140 4141 4142 4143 4144 4145 4146 4147 4148 4149
+ 4150 4151 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161 4162 4163 4164 4658 4659 4660 4661 5431
+ 5432 5433 5434
+ ICV_16 $T=364090 180630 0 0 $X=363750 $Y=180290
X1357 VSS VDD 804 4133 4134 4135 4136 4137 4138 4139 4140 4141 4142 4143 4144 4145 4146 4147 4148 4149
+ 4150 4151 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161 4162 4163 4164 4662 4663 4664 4665 5435
+ 5436 5437 5438
+ ICV_16 $T=370090 180630 0 0 $X=369750 $Y=180290
X1358 VSS VDD 804 4133 4134 4135 4136 4137 4138 4139 4140 4141 4142 4143 4144 4145 4146 4147 4148 4149
+ 4150 4151 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161 4162 4163 4164 4666 4667 4668 4669 5439
+ 5440 5441 5442
+ ICV_16 $T=376090 180630 0 0 $X=375750 $Y=180290
X1359 VSS VDD 804 4133 4134 4135 4136 4137 4138 4139 4140 4141 4142 4143 4144 4145 4146 4147 4148 4149
+ 4150 4151 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161 4162 4163 4164 4670 4671 890 889 5443
+ 5444 5445 5446
+ ICV_16 $T=382090 180630 0 0 $X=381750 $Y=180290
X1366 VSS VDD 804 4133 4134 4135 4136 4137 4138 4139 4140 4141 4142 4143 4144 4145 4146 4147 4148 4149
+ 4150 4151 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161 4162 4163 4164 4712 4713 901 900 5447
+ 5448 5449 5450
+ ICV_7 $T=340090 180630 1 180 $X=336750 $Y=180290
X1367 VSS VDD 804 4133 4134 4135 4136 4137 4138 4139 4140 4141 4142 4143 4144 4145 4146 4147 4148 4149
+ 4150 4151 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161 4162 4163 4164 4708 4709 4710 4711 5451
+ 5452 5453 5454
+ ICV_7 $T=346090 180630 1 180 $X=342750 $Y=180290
X1368 VSS VDD 804 4133 4134 4135 4136 4137 4138 4139 4140 4141 4142 4143 4144 4145 4146 4147 4148 4149
+ 4150 4151 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161 4162 4163 4164 4704 4705 4706 4707 5455
+ 5456 5457 5458
+ ICV_7 $T=352090 180630 1 180 $X=348750 $Y=180290
X1369 VSS VDD 804 4133 4134 4135 4136 4137 4138 4139 4140 4141 4142 4143 4144 4145 4146 4147 4148 4149
+ 4150 4151 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161 4162 4163 4164 4700 4701 4702 4703 5459
+ 5460 5461 5462
+ ICV_7 $T=358090 180630 1 180 $X=354750 $Y=180290
X1370 VSS VDD 804 4133 4134 4135 4136 4137 4138 4139 4140 4141 4142 4143 4144 4145 4146 4147 4148 4149
+ 4150 4151 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161 4162 4163 4164 4726 4727 904 903 5463
+ 5464 5465 5466
+ ICV_7 $T=394090 180630 1 180 $X=390750 $Y=180290
X1371 VSS VDD 804 4133 4134 4135 4136 4137 4138 4139 4140 4141 4142 4143 4144 4145 4146 4147 4148 4149
+ 4150 4151 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161 4162 4163 4164 4722 4723 4724 4725 5467
+ 5468 5469 5470
+ ICV_7 $T=400090 180630 1 180 $X=396750 $Y=180290
X1372 VSS VDD 804 4133 4134 4135 4136 4137 4138 4139 4140 4141 4142 4143 4144 4145 4146 4147 4148 4149
+ 4150 4151 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161 4162 4163 4164 4718 4719 4720 4721 5471
+ 5472 5473 5474
+ ICV_7 $T=406090 180630 1 180 $X=402750 $Y=180290
X1373 VSS VDD 804 4133 4134 4135 4136 4137 4138 4139 4140 4141 4142 4143 4144 4145 4146 4147 4148 4149
+ 4150 4151 4152 4153 4154 4155 4156 4157 4158 4159 4160 4161 4162 4163 4164 4714 4715 4716 4717 5475
+ 5476 5477 5478
+ ICV_7 $T=412090 180630 1 180 $X=408750 $Y=180290
X1382 VSS VDD 4743 4744 4745 4746 ICV_1 $T=418090 320130 0 0 $X=417750 $Y=319790
X1383 614 615 VSS VDD 4747 4748 4749 4750 ICV_2 $T=418090 176130 0 0 $X=417750 $Y=175790
X1384 614 615 VSS VDD 4751 4752 4753 4754 ICV_2 $T=418090 194130 0 0 $X=417750 $Y=193790
X1385 614 615 VSS VDD 4755 4756 4757 4758 ICV_2 $T=418090 212130 0 0 $X=417750 $Y=211790
X1386 614 615 VSS VDD 4759 4760 4761 4762 ICV_2 $T=418090 230130 0 0 $X=417750 $Y=229790
X1387 614 615 VSS VDD 4763 4764 4765 4766 ICV_2 $T=418090 248130 0 0 $X=417750 $Y=247790
X1388 614 615 VSS VDD 4767 4768 4769 4770 ICV_2 $T=418090 266130 0 0 $X=417750 $Y=265790
X1389 614 615 VSS VDD 4771 4772 4773 4774 ICV_2 $T=418090 284130 0 0 $X=417750 $Y=283790
X1390 614 615 VSS VDD 4775 4776 4777 4778 ICV_2 $T=418090 302130 0 0 $X=417750 $Y=301790
.ENDS
***************************************
