************************************************************************
* auCdl Netlist:
* 
* Library Name:  TCG_Library
* Top Cell Name: cap_pmos_06v0_b
* View Name:     schematic
* Netlisted on:  Nov 24 09:47:53 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL vdd!

*.PIN vdd!

************************************************************************
* Library Name: TCG_Library
* Cell Name:    cap_pmos_06v0_b
* View Name:    schematic
************************************************************************

.SUBCKT cap_pmos_06v0_b I1_0_0_R0_G I1_0_1_R0_G I1_0_2_R0_G I1_1_0_R0_G 
+ I1_1_1_R0_G I1_1_2_R0_G I1_2_0_R0_G I1_2_1_R0_G I1_2_2_R0_G I1_default_G vdd!
*.PININFO I1_0_0_R0_G:I I1_0_1_R0_G:I I1_0_2_R0_G:I I1_1_0_R0_G:I 
*.PININFO I1_1_1_R0_G:I I1_1_2_R0_G:I I1_2_0_R0_G:I I1_2_1_R0_G:I 
*.PININFO I1_2_2_R0_G:I I1_default_G:I vdd!:I
CI1_2_2_R0 I1_2_2_R0_G vdd! $[cap_pmos_06v0_b] m=1 l=50.000u w=50.000u
CI1_2_1_R0 I1_2_1_R0_G vdd! $[cap_pmos_06v0_b] m=1 l=50.000u w=12.350u
CI1_2_0_R0 I1_2_0_R0_G vdd! $[cap_pmos_06v0_b] m=1 l=50.000u w=1.000u
CI1_1_2_R0 I1_1_2_R0_G vdd! $[cap_pmos_06v0_b] m=1 l=12.350u w=50.000u
CI1_1_1_R0 I1_1_1_R0_G vdd! $[cap_pmos_06v0_b] m=1 l=12.350u w=12.350u
CI1_1_0_R0 I1_1_0_R0_G vdd! $[cap_pmos_06v0_b] m=1 l=12.350u w=1.000u
CI1_0_2_R0 I1_0_2_R0_G vdd! $[cap_pmos_06v0_b] m=1 l=1.000u w=50.000u
CI1_0_1_R0 I1_0_1_R0_G vdd! $[cap_pmos_06v0_b] m=1 l=1.000u w=12.350u
CI1_0_0_R0 I1_0_0_R0_G vdd! $[cap_pmos_06v0_b] m=1 l=1.000u w=1.000u
CI1_default I1_default_G vdd! $[cap_pmos_06v0_b] m=1 l=5u w=5u
.ENDS

