*Xyce Common Source Circuit
** library calling



*****************
** main netlist
*****************

Vcp c 0 dc -6
Ib 0 b -9u

xq1 c b 0 {{device}}


*****************
** Analysis
*****************
.DC Vcp 0 -3 -0.1 Ib -1u -9u -2u
.STEP TEMP {{temp}} -60 200
.print DC FORMAT=CSV file=pnp/simulated_IcVc/{{i}}_simulated_{{device}}.csv {I(Vcp)}

.include "../../../../../design.xyce"
.lib "../../../../../sm141064.xyce" bjt_typical

.end
