***************************
** pfet_03v3_t_id
***************************
* Copyright 2022 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
Vds D_tn 0 dc=-0.05
Vgs G_tn 0 dc=-6
Vbs B_tn 0 dc=0

.temp {{temp}}
 
xmp1 D_tn G_tn 0 B_tn {{device}} W = {{width}}u L = {{length}}u 

**** begin architecture code

.control
set filetype=ascii
set wr_singlescale
set wr_vecnames
dc Vgs {{vgs}} Vbs {{vbs}} 

wrdata mos_iv_regr/{{device}}/{{device}}_netlists/T{{temp}}_simulated_W{{width}}_L{{length}}.csv i(Vds) v(B_tn) v(G_tn) 
.endc

** library calling

.include "../../../design.ngspice"
.lib "../../../sm141064.ngspice" typical

**** end architecture code


.end
