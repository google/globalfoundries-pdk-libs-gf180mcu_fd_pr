*****************
** main netlist
*****************

Vcp c 0 dc -3
Vbp b 0 dc -1.2

.temp {{temp}}
.options tnom={{temp}}

xq1 c b 0 {{device}}


*****************
** Analysis
*****************

.control
set filetype=ascii

dc Vbp -0.2 -1.2 -0.01 Vcp -1 -3 -1
wrdata pnp/simulated_Ic/{{i}}_simulated_{{device}}.csv i(Vcp)
wrdata pnp/simulated_Ib/{{i}}_simulated_{{device}}.csv i(Vbp)
.endc

.include "../../../design.ngspice"
.lib "../../../sm141064.ngspice" bjt_typical

.end
