
*****************
** main netlist
*****************

Vcp c 0 dc 6
Ib 0 b 9u

.temp 25
.options tnom=25

xq1 c b 0 0 vnpn_10x10


*****************
** Analysis
*****************

.control
set filetype=ascii

dc Vcp 0 6 0.1 Ib 1u 9u 2u
print -i(Vcp)
wrdata result.csv -i(Vcp)
.endc

.include "../../../design.ngspice"
.lib "../../../sm141064.ngspice" bjt_typical

.end
