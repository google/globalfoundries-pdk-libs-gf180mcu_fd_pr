************************************************************************
* auCdl Netlist:
* 
* Library Name:  TCG_Library
* Top Cell Name: npolyf_s_dw
* View Name:     schematic
* Netlisted on:  Nov 24 09:31:45 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL gnd!

*.PIN gnd!

************************************************************************
* Library Name: TCG_Library
* Cell Name:    npolyf_s_dw
* View Name:    schematic
************************************************************************

.SUBCKT npolyf_s_dw I1_0_0_0_0_0_0_R0_MINUS I1_0_0_0_0_0_0_R0_PLUS 
+ I1_0_0_0_1_0_0_R0_MINUS I1_0_0_0_1_0_0_R0_PLUS I1_0_0_1_0_0_0_R0_MINUS 
+ I1_0_0_1_0_0_0_R0_PLUS I1_0_0_1_1_0_0_R0_MINUS I1_0_0_1_1_0_0_R0_PLUS 
+ I1_0_0_2_0_0_0_R0_MINUS I1_0_0_2_0_0_0_R0_PLUS I1_0_0_2_1_0_0_R0_MINUS 
+ I1_0_0_2_1_0_0_R0_PLUS I1_0_1_0_0_0_0_R0_MINUS I1_0_1_0_0_0_0_R0_PLUS 
+ I1_0_1_0_1_0_0_R0_MINUS I1_0_1_0_1_0_0_R0_PLUS I1_0_1_1_0_0_0_R0_MINUS 
+ I1_0_1_1_0_0_0_R0_PLUS I1_0_1_1_1_0_0_R0_MINUS I1_0_1_1_1_0_0_R0_PLUS 
+ I1_0_1_2_0_0_0_R0_MINUS I1_0_1_2_0_0_0_R0_PLUS I1_0_1_2_1_0_0_R0_MINUS 
+ I1_0_1_2_1_0_0_R0_PLUS I1_0_2_0_0_0_0_R0_MINUS I1_0_2_0_0_0_0_R0_PLUS 
+ I1_0_2_0_1_0_0_R0_MINUS I1_0_2_0_1_0_0_R0_PLUS I1_0_2_1_0_0_0_R0_MINUS 
+ I1_0_2_1_0_0_0_R0_PLUS I1_0_2_1_1_0_0_R0_MINUS I1_0_2_1_1_0_0_R0_PLUS 
+ I1_0_2_2_0_0_0_R0_MINUS I1_0_2_2_0_0_0_R0_PLUS I1_0_2_2_1_0_0_R0_MINUS 
+ I1_0_2_2_1_0_0_R0_PLUS I1_1_0_0_0_0_0_R0_MINUS I1_1_0_0_0_0_0_R0_PLUS 
+ I1_1_0_0_1_0_0_R0_MINUS I1_1_0_0_1_0_0_R0_PLUS I1_1_0_1_0_0_0_R0_MINUS 
+ I1_1_0_1_0_0_0_R0_PLUS I1_1_0_1_1_0_0_R0_MINUS I1_1_0_1_1_0_0_R0_PLUS 
+ I1_1_0_2_0_0_0_R0_MINUS I1_1_0_2_0_0_0_R0_PLUS I1_1_0_2_1_0_0_R0_MINUS 
+ I1_1_0_2_1_0_0_R0_PLUS I1_1_1_0_0_0_0_R0_MINUS I1_1_1_0_0_0_0_R0_PLUS 
+ I1_1_1_0_1_0_0_R0_MINUS I1_1_1_0_1_0_0_R0_PLUS I1_1_1_1_0_0_0_R0_MINUS 
+ I1_1_1_1_0_0_0_R0_PLUS I1_1_1_1_1_0_0_R0_MINUS I1_1_1_1_1_0_0_R0_PLUS 
+ I1_1_1_2_0_0_0_R0_MINUS I1_1_1_2_0_0_0_R0_PLUS I1_1_1_2_1_0_0_R0_MINUS 
+ I1_1_1_2_1_0_0_R0_PLUS I1_1_2_0_0_0_0_R0_MINUS I1_1_2_0_0_0_0_R0_PLUS 
+ I1_1_2_0_1_0_0_R0_MINUS I1_1_2_0_1_0_0_R0_PLUS I1_1_2_1_0_0_0_R0_MINUS 
+ I1_1_2_1_0_0_0_R0_PLUS I1_1_2_1_1_0_0_R0_MINUS I1_1_2_1_1_0_0_R0_PLUS 
+ I1_1_2_2_0_0_0_R0_MINUS I1_1_2_2_0_0_0_R0_PLUS I1_1_2_2_1_0_0_R0_MINUS 
+ I1_1_2_2_1_0_0_R0_PLUS I1_2_0_0_0_0_0_R0_MINUS I1_2_0_0_0_0_0_R0_PLUS 
+ I1_2_0_0_1_0_0_R0_MINUS I1_2_0_0_1_0_0_R0_PLUS I1_2_0_1_0_0_0_R0_MINUS 
+ I1_2_0_1_0_0_0_R0_PLUS I1_2_0_1_1_0_0_R0_MINUS I1_2_0_1_1_0_0_R0_PLUS 
+ I1_2_0_2_0_0_0_R0_MINUS I1_2_0_2_0_0_0_R0_PLUS I1_2_0_2_1_0_0_R0_MINUS 
+ I1_2_0_2_1_0_0_R0_PLUS I1_2_1_0_0_0_0_R0_MINUS I1_2_1_0_0_0_0_R0_PLUS 
+ I1_2_1_0_1_0_0_R0_MINUS I1_2_1_0_1_0_0_R0_PLUS I1_2_1_1_0_0_0_R0_MINUS 
+ I1_2_1_1_0_0_0_R0_PLUS I1_2_1_1_1_0_0_R0_MINUS I1_2_1_1_1_0_0_R0_PLUS 
+ I1_2_1_2_0_0_0_R0_MINUS I1_2_1_2_0_0_0_R0_PLUS I1_2_1_2_1_0_0_R0_MINUS 
+ I1_2_1_2_1_0_0_R0_PLUS I1_2_2_0_0_0_0_R0_MINUS I1_2_2_0_0_0_0_R0_PLUS 
+ I1_2_2_0_1_0_0_R0_MINUS I1_2_2_0_1_0_0_R0_PLUS I1_2_2_1_0_0_0_R0_MINUS 
+ I1_2_2_1_0_0_0_R0_PLUS I1_2_2_1_1_0_0_R0_MINUS I1_2_2_1_1_0_0_R0_PLUS 
+ I1_2_2_2_0_0_0_R0_MINUS I1_2_2_2_0_0_0_R0_PLUS I1_2_2_2_1_0_0_R0_MINUS 
+ I1_2_2_2_1_0_0_R0_PLUS I1_default_MINUS I1_default_PLUS gnd!
*.PININFO I1_0_0_0_0_0_0_R0_MINUS:I I1_0_0_0_0_0_0_R0_PLUS:I 
*.PININFO I1_0_0_0_1_0_0_R0_MINUS:I I1_0_0_0_1_0_0_R0_PLUS:I 
*.PININFO I1_0_0_1_0_0_0_R0_MINUS:I I1_0_0_1_0_0_0_R0_PLUS:I 
*.PININFO I1_0_0_1_1_0_0_R0_MINUS:I I1_0_0_1_1_0_0_R0_PLUS:I 
*.PININFO I1_0_0_2_0_0_0_R0_MINUS:I I1_0_0_2_0_0_0_R0_PLUS:I 
*.PININFO I1_0_0_2_1_0_0_R0_MINUS:I I1_0_0_2_1_0_0_R0_PLUS:I 
*.PININFO I1_0_1_0_0_0_0_R0_MINUS:I I1_0_1_0_0_0_0_R0_PLUS:I 
*.PININFO I1_0_1_0_1_0_0_R0_MINUS:I I1_0_1_0_1_0_0_R0_PLUS:I 
*.PININFO I1_0_1_1_0_0_0_R0_MINUS:I I1_0_1_1_0_0_0_R0_PLUS:I 
*.PININFO I1_0_1_1_1_0_0_R0_MINUS:I I1_0_1_1_1_0_0_R0_PLUS:I 
*.PININFO I1_0_1_2_0_0_0_R0_MINUS:I I1_0_1_2_0_0_0_R0_PLUS:I 
*.PININFO I1_0_1_2_1_0_0_R0_MINUS:I I1_0_1_2_1_0_0_R0_PLUS:I 
*.PININFO I1_0_2_0_0_0_0_R0_MINUS:I I1_0_2_0_0_0_0_R0_PLUS:I 
*.PININFO I1_0_2_0_1_0_0_R0_MINUS:I I1_0_2_0_1_0_0_R0_PLUS:I 
*.PININFO I1_0_2_1_0_0_0_R0_MINUS:I I1_0_2_1_0_0_0_R0_PLUS:I 
*.PININFO I1_0_2_1_1_0_0_R0_MINUS:I I1_0_2_1_1_0_0_R0_PLUS:I 
*.PININFO I1_0_2_2_0_0_0_R0_MINUS:I I1_0_2_2_0_0_0_R0_PLUS:I 
*.PININFO I1_0_2_2_1_0_0_R0_MINUS:I I1_0_2_2_1_0_0_R0_PLUS:I 
*.PININFO I1_1_0_0_0_0_0_R0_MINUS:I I1_1_0_0_0_0_0_R0_PLUS:I 
*.PININFO I1_1_0_0_1_0_0_R0_MINUS:I I1_1_0_0_1_0_0_R0_PLUS:I 
*.PININFO I1_1_0_1_0_0_0_R0_MINUS:I I1_1_0_1_0_0_0_R0_PLUS:I 
*.PININFO I1_1_0_1_1_0_0_R0_MINUS:I I1_1_0_1_1_0_0_R0_PLUS:I 
*.PININFO I1_1_0_2_0_0_0_R0_MINUS:I I1_1_0_2_0_0_0_R0_PLUS:I 
*.PININFO I1_1_0_2_1_0_0_R0_MINUS:I I1_1_0_2_1_0_0_R0_PLUS:I 
*.PININFO I1_1_1_0_0_0_0_R0_MINUS:I I1_1_1_0_0_0_0_R0_PLUS:I 
*.PININFO I1_1_1_0_1_0_0_R0_MINUS:I I1_1_1_0_1_0_0_R0_PLUS:I 
*.PININFO I1_1_1_1_0_0_0_R0_MINUS:I I1_1_1_1_0_0_0_R0_PLUS:I 
*.PININFO I1_1_1_1_1_0_0_R0_MINUS:I I1_1_1_1_1_0_0_R0_PLUS:I 
*.PININFO I1_1_1_2_0_0_0_R0_MINUS:I I1_1_1_2_0_0_0_R0_PLUS:I 
*.PININFO I1_1_1_2_1_0_0_R0_MINUS:I I1_1_1_2_1_0_0_R0_PLUS:I 
*.PININFO I1_1_2_0_0_0_0_R0_MINUS:I I1_1_2_0_0_0_0_R0_PLUS:I 
*.PININFO I1_1_2_0_1_0_0_R0_MINUS:I I1_1_2_0_1_0_0_R0_PLUS:I 
*.PININFO I1_1_2_1_0_0_0_R0_MINUS:I I1_1_2_1_0_0_0_R0_PLUS:I 
*.PININFO I1_1_2_1_1_0_0_R0_MINUS:I I1_1_2_1_1_0_0_R0_PLUS:I 
*.PININFO I1_1_2_2_0_0_0_R0_MINUS:I I1_1_2_2_0_0_0_R0_PLUS:I 
*.PININFO I1_1_2_2_1_0_0_R0_MINUS:I I1_1_2_2_1_0_0_R0_PLUS:I 
*.PININFO I1_2_0_0_0_0_0_R0_MINUS:I I1_2_0_0_0_0_0_R0_PLUS:I 
*.PININFO I1_2_0_0_1_0_0_R0_MINUS:I I1_2_0_0_1_0_0_R0_PLUS:I 
*.PININFO I1_2_0_1_0_0_0_R0_MINUS:I I1_2_0_1_0_0_0_R0_PLUS:I 
*.PININFO I1_2_0_1_1_0_0_R0_MINUS:I I1_2_0_1_1_0_0_R0_PLUS:I 
*.PININFO I1_2_0_2_0_0_0_R0_MINUS:I I1_2_0_2_0_0_0_R0_PLUS:I 
*.PININFO I1_2_0_2_1_0_0_R0_MINUS:I I1_2_0_2_1_0_0_R0_PLUS:I 
*.PININFO I1_2_1_0_0_0_0_R0_MINUS:I I1_2_1_0_0_0_0_R0_PLUS:I 
*.PININFO I1_2_1_0_1_0_0_R0_MINUS:I I1_2_1_0_1_0_0_R0_PLUS:I 
*.PININFO I1_2_1_1_0_0_0_R0_MINUS:I I1_2_1_1_0_0_0_R0_PLUS:I 
*.PININFO I1_2_1_1_1_0_0_R0_MINUS:I I1_2_1_1_1_0_0_R0_PLUS:I 
*.PININFO I1_2_1_2_0_0_0_R0_MINUS:I I1_2_1_2_0_0_0_R0_PLUS:I 
*.PININFO I1_2_1_2_1_0_0_R0_MINUS:I I1_2_1_2_1_0_0_R0_PLUS:I 
*.PININFO I1_2_2_0_0_0_0_R0_MINUS:I I1_2_2_0_0_0_0_R0_PLUS:I 
*.PININFO I1_2_2_0_1_0_0_R0_MINUS:I I1_2_2_0_1_0_0_R0_PLUS:I 
*.PININFO I1_2_2_1_0_0_0_R0_MINUS:I I1_2_2_1_0_0_0_R0_PLUS:I 
*.PININFO I1_2_2_1_1_0_0_R0_MINUS:I I1_2_2_1_1_0_0_R0_PLUS:I 
*.PININFO I1_2_2_2_0_0_0_R0_MINUS:I I1_2_2_2_0_0_0_R0_PLUS:I 
*.PININFO I1_2_2_2_1_0_0_R0_MINUS:I I1_2_2_2_1_0_0_R0_PLUS:I 
*.PININFO I1_default_MINUS:I I1_default_PLUS:I gnd!:I
RI1_2_2_2_1_0_0_R0 I1_2_2_2_1_0_0_R0_PLUS I1_2_2_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=8.0 l=50u w=50u r=7.02182 par=8.0 s=1
RI1_2_2_2_0_0_0_R0 I1_2_2_2_0_0_0_R0_PLUS I1_2_2_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=50u w=50u r=7.02182 par=1.0 s=8
RI1_2_2_1_1_0_0_R0 I1_2_2_1_1_0_0_R0_PLUS I1_2_2_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=3.0 l=50u w=50u r=7.02182 par=3.0 s=1
RI1_2_2_1_0_0_0_R0 I1_2_2_1_0_0_0_R0_PLUS I1_2_2_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=50u w=50u r=7.02182 par=1.0 s=3
RI1_2_2_0_1_0_0_R0 I1_2_2_0_1_0_0_R0_PLUS I1_2_2_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=50u w=50u r=7.02182 par=1.0 s=1
RI1_2_2_0_0_0_0_R0 I1_2_2_0_0_0_0_R0_PLUS I1_2_2_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=50u w=50u r=7.02182 par=1.0 s=1
RI1_2_1_2_1_0_0_R0 I1_2_1_2_1_0_0_R0_PLUS I1_2_1_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=8.0 l=7.6u w=50u r=1.25392 par=8.0 s=1
RI1_2_1_2_0_0_0_R0 I1_2_1_2_0_0_0_R0_PLUS I1_2_1_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=7.6u w=50u r=1.25392 par=1.0 s=8
RI1_2_1_1_1_0_0_R0 I1_2_1_1_1_0_0_R0_PLUS I1_2_1_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=3.0 l=7.6u w=50u r=1.25392 par=3.0 s=1
RI1_2_1_1_0_0_0_R0 I1_2_1_1_0_0_0_R0_PLUS I1_2_1_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=7.6u w=50u r=1.25392 par=1.0 s=3
RI1_2_1_0_1_0_0_R0 I1_2_1_0_1_0_0_R0_PLUS I1_2_1_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=7.6u w=50u r=1.25392 par=1.0 s=1
RI1_2_1_0_0_0_0_R0 I1_2_1_0_0_0_0_R0_PLUS I1_2_1_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=7.6u w=50u r=1.25392 par=1.0 s=1
RI1_2_0_2_1_0_0_R0 I1_2_0_2_1_0_0_R0_PLUS I1_2_0_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=8.0 l=1.6u w=50u r=437.71m par=8.0 s=1
RI1_2_0_2_0_0_0_R0 I1_2_0_2_0_0_0_R0_PLUS I1_2_0_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=1.6u w=50u r=437.71m par=1.0 s=8
RI1_2_0_1_1_0_0_R0 I1_2_0_1_1_0_0_R0_PLUS I1_2_0_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=3.0 l=1.6u w=50u r=437.71m par=3.0 s=1
RI1_2_0_1_0_0_0_R0 I1_2_0_1_0_0_0_R0_PLUS I1_2_0_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=1.6u w=50u r=437.71m par=1.0 s=3
RI1_2_0_0_1_0_0_R0 I1_2_0_0_1_0_0_R0_PLUS I1_2_0_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=1.6u w=50u r=437.71m par=1.0 s=1
RI1_2_0_0_0_0_0_R0 I1_2_0_0_0_0_0_R0_PLUS I1_2_0_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=1.6u w=50u r=437.71m par=1.0 s=1
RI1_1_2_2_1_0_0_R0 I1_1_2_2_1_0_0_R0_PLUS I1_1_2_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=8.0 l=50u w=3.62u r=97.3107 par=8.0 s=1
RI1_1_2_2_0_0_0_R0 I1_1_2_2_0_0_0_R0_PLUS I1_1_2_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=50u w=3.62u r=97.3107 par=1.0 s=8
RI1_1_2_1_1_0_0_R0 I1_1_2_1_1_0_0_R0_PLUS I1_1_2_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=3.0 l=50u w=3.62u r=97.3107 par=3.0 s=1
RI1_1_2_1_0_0_0_R0 I1_1_2_1_0_0_0_R0_PLUS I1_1_2_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=50u w=3.62u r=97.3107 par=1.0 s=3
RI1_1_2_0_1_0_0_R0 I1_1_2_0_1_0_0_R0_PLUS I1_1_2_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=50u w=3.62u r=97.3107 par=1.0 s=1
RI1_1_2_0_0_0_0_R0 I1_1_2_0_0_0_0_R0_PLUS I1_1_2_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=50u w=3.62u r=97.3107 par=1.0 s=1
RI1_1_1_2_1_0_0_R0 I1_1_1_2_1_0_0_R0_PLUS I1_1_1_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=8.0 l=7.6u w=3.62u r=17.3773 par=8.0 s=1
RI1_1_1_2_0_0_0_R0 I1_1_1_2_0_0_0_R0_PLUS I1_1_1_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=7.6u w=3.62u r=17.3773 par=1.0 s=8
RI1_1_1_1_1_0_0_R0 I1_1_1_1_1_0_0_R0_PLUS I1_1_1_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=3.0 l=7.6u w=3.62u r=17.3773 par=3.0 s=1
RI1_1_1_1_0_0_0_R0 I1_1_1_1_0_0_0_R0_PLUS I1_1_1_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=7.6u w=3.62u r=17.3773 par=1.0 s=3
RI1_1_1_0_1_0_0_R0 I1_1_1_0_1_0_0_R0_PLUS I1_1_1_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=7.6u w=3.62u r=17.3773 par=1.0 s=1
RI1_1_1_0_0_0_0_R0 I1_1_1_0_0_0_0_R0_PLUS I1_1_1_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=7.6u w=3.62u r=17.3773 par=1.0 s=1
RI1_1_0_2_1_0_0_R0 I1_1_0_2_1_0_0_R0_PLUS I1_1_0_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=8.0 l=1.6u w=3.62u r=6.06593 par=8.0 s=1
RI1_1_0_2_0_0_0_R0 I1_1_0_2_0_0_0_R0_PLUS I1_1_0_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=1.6u w=3.62u r=6.06593 par=1.0 s=8
RI1_1_0_1_1_0_0_R0 I1_1_0_1_1_0_0_R0_PLUS I1_1_0_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=3.0 l=1.6u w=3.62u r=6.06593 par=3.0 s=1
RI1_1_0_1_0_0_0_R0 I1_1_0_1_0_0_0_R0_PLUS I1_1_0_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=1.6u w=3.62u r=6.06593 par=1.0 s=3
RI1_1_0_0_1_0_0_R0 I1_1_0_0_1_0_0_R0_PLUS I1_1_0_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=1.6u w=3.62u r=6.06593 par=1.0 s=1
RI1_1_0_0_0_0_0_R0 I1_1_0_0_0_0_0_R0_PLUS I1_1_0_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=1.6u w=3.62u r=6.06593 par=1.0 s=1
RI1_0_2_2_1_0_0_R0 I1_0_2_2_1_0_0_R0_PLUS I1_0_2_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=8.0 l=50u w=800n r=445.997 par=8.0 s=1
RI1_0_2_2_0_0_0_R0 I1_0_2_2_0_0_0_R0_PLUS I1_0_2_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=50u w=800n r=445.997 par=1.0 s=8
RI1_0_2_1_1_0_0_R0 I1_0_2_1_1_0_0_R0_PLUS I1_0_2_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=3.0 l=50u w=800n r=445.997 par=3.0 s=1
RI1_0_2_1_0_0_0_R0 I1_0_2_1_0_0_0_R0_PLUS I1_0_2_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=50u w=800n r=445.997 par=1.0 s=3
RI1_0_2_0_1_0_0_R0 I1_0_2_0_1_0_0_R0_PLUS I1_0_2_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=50u w=800n r=445.997 par=1.0 s=1
RI1_0_2_0_0_0_0_R0 I1_0_2_0_0_0_0_R0_PLUS I1_0_2_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=50u w=800n r=445.997 par=1.0 s=1
RI1_0_1_2_1_0_0_R0 I1_0_1_2_1_0_0_R0_PLUS I1_0_1_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=8.0 l=7.6u w=800n r=79.644 par=8.0 s=1
RI1_0_1_2_0_0_0_R0 I1_0_1_2_0_0_0_R0_PLUS I1_0_1_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=7.6u w=800n r=79.644 par=1.0 s=8
RI1_0_1_1_1_0_0_R0 I1_0_1_1_1_0_0_R0_PLUS I1_0_1_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=3.0 l=7.6u w=800n r=79.644 par=3.0 s=1
RI1_0_1_1_0_0_0_R0 I1_0_1_1_0_0_0_R0_PLUS I1_0_1_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=7.6u w=800n r=79.644 par=1.0 s=3
RI1_0_1_0_1_0_0_R0 I1_0_1_0_1_0_0_R0_PLUS I1_0_1_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=7.6u w=800n r=79.644 par=1.0 s=1
RI1_0_1_0_0_0_0_R0 I1_0_1_0_0_0_0_R0_PLUS I1_0_1_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=7.6u w=800n r=79.644 par=1.0 s=1
RI1_0_0_2_1_0_0_R0 I1_0_0_2_1_0_0_R0_PLUS I1_0_0_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=8.0 l=1.6u w=800n r=27.8015 par=8.0 s=1
RI1_0_0_2_0_0_0_R0 I1_0_0_2_0_0_0_R0_PLUS I1_0_0_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=1.6u w=800n r=27.8015 par=1.0 s=8
RI1_0_0_1_1_0_0_R0 I1_0_0_1_1_0_0_R0_PLUS I1_0_0_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=3.0 l=1.6u w=800n r=27.8015 par=3.0 s=1
RI1_0_0_1_0_0_0_R0 I1_0_0_1_0_0_0_R0_PLUS I1_0_0_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=1.6u w=800n r=27.8015 par=1.0 s=3
RI1_0_0_0_1_0_0_R0 I1_0_0_0_1_0_0_R0_PLUS I1_0_0_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=1.6u w=800n r=27.8015 par=1.0 s=1
RI1_0_0_0_0_0_0_R0 I1_0_0_0_0_0_0_R0_PLUS I1_0_0_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[npolyf_s_dw] m=1.0 l=1.6u w=800n r=27.8015 par=1.0 s=1
RI1_default I1_default_PLUS I1_default_MINUS $SUB=gnd! $[npolyf_s_dw] m=1.0 
+ l=1.6u w=800.0n r=27.8015 par=1.0 s=1
.ENDS

