*****************
** BJT-iv netlist
*****************
* Copyright 2023 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

Vcp c 0 dc=6
Ib f b 9u
Vbb 0 f dc=0

.temp {{temp}}

xq {{terminals}} {{device}}

*****************
** Analysis
*****************
.control
set filetype=ascii
set wr_singlescale
set wr_vecnames

dc {{sweep}}

let vcp = v(c)
let ibp = i(Vbb)
let ic = -i(Vcp)

wrdata {{result_path}} ibp vcp ic 
.endc

** library calling

.include {{model_design_path}}
.lib {{model_card_path}} {{corner}}

**** end architecture code

.end
