**************************
** res
**************************
* Copyright 2022 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

Vin top GND {{voltage}}
XR1 top {{terminals}} {{device}} r_width={{width}}u r_length={{length}}u m=1

.temp {{temp}}
.options tnom={{temp}}

.control
op
let ires=-1*vin#branch
let res={{voltage}}/ires
print res
.endc

** library calling

.include "../../../design.ngspice"
.lib "../../../sm141064.ngspice" res_{{corner}}

.GLOBAL GND
.end