***************************
** cap
***************************
* Copyright 2022 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
.options noacct

Ich 0 p dc 10u

.temp 25
.options tnom=25
      
xcn p 0 cap_nmos_03v3_b c_length=1.0u c_width=50.0u

.ic v(p)=0.0
.tran 10ns 100us

* .print tran v(p) cj=par('10.0e-6  * time / v(p)')

.meas tran CV FIND par('(10.0e-6  * time / v(p))*1.0e15') AT=100us

** library calling

.include "../../../design.ngspice"
.lib "../../../sm141064.ngspice" moscap_ff
.end
