*Xyce Common Source Circuit
** library calling



*****************
** main netlist
*****************
Vds D_tn 0 dc -3.3
Vgs G_tn 0 dc -3.3


xmn1 D_tn G_tn 0 0 pmos_3p3_sab W={{width}}u L={{length}}u ad={{AD}}u pd={{PD}}u as={{AS}}u ps={{PS}}u



*****************
** Analysis
*****************
.DC Vds 0 -3.3 -0.05 Vgs -0.8 -3.3 -0.5
.STEP TEMP {{temp}} -60 200
.print DC FORMAT=CSV file=pmos_3p3_sab_iv/simulated_Rds/{{i}}_simulated_W{{width}}_L{{length}}.csv {1/N(xmn1:m0:gds)}

.include "../../../../../design.xyce"
.lib "../../../../../sm141064.xyce" typical

.end