**************************
** res
**************************
* Copyright 2022 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

Vn n 0 DC {{sign}}3.3

.temp {{temp}}
.options tnom={{temp}}
      
r1 n p 1M
xrn p 0 {{device}} r_width={{width}}u r_length={{length}}u


.print dc Rs=par('(1M*V(p)/(V(n)-V(p)))/{{length}}u*{{width}}u')


.control
set filetype=ascii
set appendwrite

DC Vn {{sign}}3.3 {{sign}}3.3 0.1
wrdata {{device}}_r_{{corner}}_temp/simulated_r/{{i}}_simulated_w{{width}}_l{{length}}.csv Rs 

.endc

** library calling

.include "../../../design.ngspice"
.lib "../../../sm141064.ngspice" res_{{corner}}

.end
