**********************
** DIODE-IV netlist **
**********************
* Copyright 2023 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
Vn n 0 dc=1

.temp {{temp}}
.options GMIN=1.0e-16 ABSTOL=1e-15

dn n 0 {{device}} AREA = {{area}}p PJ = {{perim}}u 

**** begin architecture code

.control
set filetype=ascii
set wr_singlescale
set wr_vecnames

dc {{sweep}}

let In = abs(i(Vn))
let Vn = V(n)

wrdata {{result_path}} Vn In
.endc

** library calling

.include {{model_design_path}}
.lib {{model_card_path}} {{corner}}

**** end architecture code

.end
