*Xyce Common Source Circuit
** library calling



*****************
** main netlist
*****************
.param volt = -3.0
V1 in 0 dc {volt} ac 1
*Iopen open 0 0

R1 in out 1G
xq1 0 out 0 0 vnpn_10x10

.meas AC freq when Vdb(out)=-3 PRECISION=15

*****************
** Analysis
*****************
.ac dec 10 1 10G
.STEP volt 0 -3.0 -0.1
.STEP TEMP 25 -60 200

.include "../../../../design.xyce"
.lib "../../../../sm141064.xyce" bjt_typical

.end
