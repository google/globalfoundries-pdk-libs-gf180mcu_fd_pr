************************************************************************
* auCdl Netlist:
* 
* Library Name:  TCG_Library
* Top Cell Name: tm6k
* View Name:     schematic
* Netlisted on:  Nov 24 10:55:47 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: TCG_Library
* Cell Name:    tm6k
* View Name:    schematic
************************************************************************

.SUBCKT tm6k
*.PININFO
RI1_2_2_R0 net1 net2 $[tm6k] $W=50u $L=50u m=1 r=60m par=1 dtemp=0
RI1_2_1_R0 net3 net4 $[tm6k] $W=50u $L=13.5u m=1 r=16.2m par=1 dtemp=0
RI1_2_0_R0 net5 net6 $[tm6k] $W=50u $L=360n m=1 r=432u par=1 dtemp=0
RI1_1_2_R0 net7 net8 $[tm6k] $W=13.5u $L=50u m=1 r=222.222m par=1 dtemp=0
RI1_1_1_R0 net9 net10 $[tm6k] $W=13.5u $L=13.5u m=1 r=60m par=1 dtemp=0
RI1_1_0_R0 net11 net12 $[tm6k] $W=13.5u $L=360n m=1 r=1.6m par=1 dtemp=0
RI1_0_2_R0 net13 net14 $[tm6k] $W=360n $L=50u m=1 r=8.33333 par=1 dtemp=0
RI1_0_1_R0 net15 net16 $[tm6k] $W=360n $L=13.5u m=1 r=2.25 par=1 dtemp=0
RI1_0_0_R0 net17 net18 $[tm6k] $W=360n $L=360n m=1 r=60m par=1 dtemp=0
RI1_default net19 net20 $[tm6k] $W=360.00n $L=360.00n m=1 r=60.00m par=1 
+ dtemp=0
.ENDS

