*Xyce Common Source Circuit
** library calling

* .OPTIONS DEVICE TEMP=-40

*****************
** main netlist
*****************
Vds D_tn 0 dc 3.3
Vgs G_tn 0 dc 3.3


xmn1 D_tn G_tn 0 0 nmos_6p0_nat W={{width}}u L={{length}}u ad={{AD}}u pd={{PD}}u as={{AS}}u ps={{PS}}u

*****************
** Analysis
*****************
.DC Vds 0 6.6 0.05 Vgs 0.25 6 1.15
.STEP TEMP {{temp}} -60 200
.print DC FORMAT=CSV file=nmos_6p0_nat_iv/simulated_Id/{{i}}_simulated_W{{width}}_L{{length}}.csv {-I(Vds)}

.include "../../../../../design.xyce"
.lib "../../../../../sm141064.xyce" typical

.end