************************************************************************
* auCdl Netlist:
* 
* Library Name:  TCG_Library
* Top Cell Name: mim_2p0fF_tm
* View Name:     schematic
* Netlisted on:  Nov 24 11:32:36 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: TCG_Library
* Cell Name:    mim_2p0fF_tm
* View Name:    schematic
************************************************************************

.SUBCKT mim_2p0fF_tm I1_0_0_R0_BOT I1_0_0_R0_TOP I1_0_1_R0_BOT I1_0_1_R0_TOP 
+ I1_0_2_R0_BOT I1_0_2_R0_TOP I1_1_0_R0_BOT I1_1_0_R0_TOP I1_1_1_R0_BOT 
+ I1_1_1_R0_TOP I1_1_2_R0_BOT I1_1_2_R0_TOP I1_2_0_R0_BOT I1_2_0_R0_TOP 
+ I1_2_1_R0_BOT I1_2_1_R0_TOP I1_2_2_R0_BOT I1_2_2_R0_TOP I1_default_BOT 
+ I1_default_TOP
*.PININFO I1_0_0_R0_BOT:I I1_0_0_R0_TOP:I I1_0_1_R0_BOT:I I1_0_1_R0_TOP:I 
*.PININFO I1_0_2_R0_BOT:I I1_0_2_R0_TOP:I I1_1_0_R0_BOT:I I1_1_0_R0_TOP:I 
*.PININFO I1_1_1_R0_BOT:I I1_1_1_R0_TOP:I I1_1_2_R0_BOT:I I1_1_2_R0_TOP:I 
*.PININFO I1_2_0_R0_BOT:I I1_2_0_R0_TOP:I I1_2_1_R0_BOT:I I1_2_1_R0_TOP:I 
*.PININFO I1_2_2_R0_BOT:I I1_2_2_R0_TOP:I I1_default_BOT:I I1_default_TOP:I
CI1_2_2_R0 I1_2_2_R0_TOP I1_2_2_R0_BOT $[mim_single_2p0fF] M=1 l=100.000u 
+ w=100.000u c=19.99532p
CI1_2_1_R0 I1_2_1_R0_TOP I1_2_1_R0_BOT $[mim_single_2p0fF] M=1 l=100.000u 
+ w=12.340u c=2.50920124p
CI1_2_0_R0 I1_2_0_R0_TOP I1_2_0_R0_BOT $[mim_single_2p0fF] M=1 l=100.000u 
+ w=5.000u c=1.045043p
CI1_1_2_R0 I1_1_2_R0_TOP I1_1_2_R0_BOT $[mim_single_2p0fF] M=1 l=12.340u 
+ w=100.000u c=2.50920124p
CI1_1_1_R0 I1_1_1_R0_TOP I1_1_1_R0_BOT $[mim_single_2p0fF] M=1 l=12.340u 
+ w=12.340u c=0.31479093p
CI1_1_0_R0 I1_1_0_R0_TOP I1_1_0_R0_BOT $[mim_single_2p0fF] M=1 l=12.340u 
+ w=5.000u c=0.13104724p
CI1_0_2_R0 I1_0_2_R0_TOP I1_0_2_R0_BOT $[mim_single_2p0fF] M=1 l=5.000u 
+ w=100.000u c=1.045043p
CI1_0_1_R0 I1_0_1_R0_TOP I1_0_1_R0_BOT $[mim_single_2p0fF] M=1 l=5.000u 
+ w=12.340u c=0.13104724p
CI1_0_0_R0 I1_0_0_R0_TOP I1_0_0_R0_BOT $[mim_single_2p0fF] M=1 l=5.000u 
+ w=5.000u c=0.054516p
CI1_default I1_default_TOP I1_default_BOT $[mim_single_2p0fF] M=1 l=5u w=5u 
+ c=0.054516p
.ENDS

