* ***************************
* ** pfet_03v3_t_Rds
* ***************************
* * Copyright 2023 Efabless Corporation
* *
* * Licensed under the Apache License, Version 2.0 (the "License");
* * you may not use this file except in compliance with the License.
* * You may obtain a copy of the License at
* *
* *      http://www.apache.org/licenses/LICENSE-2.0
* *
* * Unless required by applicable law or agreed to in writing, software
* * distributed under the License is distributed on an "AS IS" BASIS,
* * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* * See the License for the specific language governing permissions and
* * limitations under the License.

vds D_tn 0 dc={{vds_val}}
vgs G_tn 0 dc=-3.3
Vbs B_tn 0 dc={{vbs_val}}

.temp {{temp}} 

xmp1 D_tn G_tn 0 0 {{device}} W = {{width}}u L = {{length}}u

**** begin architecture code

.control
set filetype=ascii
set wr_singlescale
set wr_vecnames
dc {{sweeps}}

** Get all voltages and currrent
let vds = v(D_tn)
let vgs = v(G_tn)
let vbs = v(B_tn)
let rds = 1/deriv(-i(Vds))

wrdata mos_iv_regr/{{device}}/{{device}}_netlists/simulated_w{{width}}_l{{length}}_t{{temp}}_{{const_var}}{{const_var_val}}_{{meas_out_result}}.csv vds vgs vbs rds
.endc

** library calling

.include "../../../design.ngspice"
.lib "../../../sm141064.ngspice" typical

**** end architecture code

.end
