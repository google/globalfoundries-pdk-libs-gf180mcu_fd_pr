************************************************************************
* auCdl Netlist:
* 
* Library Name:  TCG_Library
* Top Cell Name: nplus_s_dw
* View Name:     schematic
* Netlisted on:  Nov 24 09:25:53 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL gnd!

*.PIN gnd!

************************************************************************
* Library Name: TCG_Library
* Cell Name:    nplus_s_dw
* View Name:    schematic
************************************************************************

.SUBCKT nplus_s_dw I1_0_0_0_0_0_0_R0_MINUS I1_0_0_0_0_0_0_R0_PLUS 
+ I1_0_0_0_1_0_0_R0_MINUS I1_0_0_0_1_0_0_R0_PLUS I1_0_0_1_0_0_0_R0_MINUS 
+ I1_0_0_1_0_0_0_R0_PLUS I1_0_0_1_1_0_0_R0_MINUS I1_0_0_1_1_0_0_R0_PLUS 
+ I1_0_0_2_0_0_0_R0_MINUS I1_0_0_2_0_0_0_R0_PLUS I1_0_0_2_1_0_0_R0_MINUS 
+ I1_0_0_2_1_0_0_R0_PLUS I1_0_1_0_0_0_0_R0_MINUS I1_0_1_0_0_0_0_R0_PLUS 
+ I1_0_1_0_1_0_0_R0_MINUS I1_0_1_0_1_0_0_R0_PLUS I1_0_1_1_0_0_0_R0_MINUS 
+ I1_0_1_1_0_0_0_R0_PLUS I1_0_1_1_1_0_0_R0_MINUS I1_0_1_1_1_0_0_R0_PLUS 
+ I1_0_1_2_0_0_0_R0_MINUS I1_0_1_2_0_0_0_R0_PLUS I1_0_1_2_1_0_0_R0_MINUS 
+ I1_0_1_2_1_0_0_R0_PLUS I1_0_2_0_0_0_0_R0_MINUS I1_0_2_0_0_0_0_R0_PLUS 
+ I1_0_2_0_1_0_0_R0_MINUS I1_0_2_0_1_0_0_R0_PLUS I1_0_2_1_0_0_0_R0_MINUS 
+ I1_0_2_1_0_0_0_R0_PLUS I1_0_2_1_1_0_0_R0_MINUS I1_0_2_1_1_0_0_R0_PLUS 
+ I1_0_2_2_0_0_0_R0_MINUS I1_0_2_2_0_0_0_R0_PLUS I1_0_2_2_1_0_0_R0_MINUS 
+ I1_0_2_2_1_0_0_R0_PLUS I1_1_0_0_0_0_0_R0_MINUS I1_1_0_0_0_0_0_R0_PLUS 
+ I1_1_0_0_1_0_0_R0_MINUS I1_1_0_0_1_0_0_R0_PLUS I1_1_0_1_0_0_0_R0_MINUS 
+ I1_1_0_1_0_0_0_R0_PLUS I1_1_0_1_1_0_0_R0_MINUS I1_1_0_1_1_0_0_R0_PLUS 
+ I1_1_0_2_0_0_0_R0_MINUS I1_1_0_2_0_0_0_R0_PLUS I1_1_0_2_1_0_0_R0_MINUS 
+ I1_1_0_2_1_0_0_R0_PLUS I1_1_1_0_0_0_0_R0_MINUS I1_1_1_0_0_0_0_R0_PLUS 
+ I1_1_1_0_1_0_0_R0_MINUS I1_1_1_0_1_0_0_R0_PLUS I1_1_1_1_0_0_0_R0_MINUS 
+ I1_1_1_1_0_0_0_R0_PLUS I1_1_1_1_1_0_0_R0_MINUS I1_1_1_1_1_0_0_R0_PLUS 
+ I1_1_1_2_0_0_0_R0_MINUS I1_1_1_2_0_0_0_R0_PLUS I1_1_1_2_1_0_0_R0_MINUS 
+ I1_1_1_2_1_0_0_R0_PLUS I1_1_2_0_0_0_0_R0_MINUS I1_1_2_0_0_0_0_R0_PLUS 
+ I1_1_2_0_1_0_0_R0_MINUS I1_1_2_0_1_0_0_R0_PLUS I1_1_2_1_0_0_0_R0_MINUS 
+ I1_1_2_1_0_0_0_R0_PLUS I1_1_2_1_1_0_0_R0_MINUS I1_1_2_1_1_0_0_R0_PLUS 
+ I1_1_2_2_0_0_0_R0_MINUS I1_1_2_2_0_0_0_R0_PLUS I1_1_2_2_1_0_0_R0_MINUS 
+ I1_1_2_2_1_0_0_R0_PLUS I1_2_0_0_0_0_0_R0_MINUS I1_2_0_0_0_0_0_R0_PLUS 
+ I1_2_0_0_1_0_0_R0_MINUS I1_2_0_0_1_0_0_R0_PLUS I1_2_0_1_0_0_0_R0_MINUS 
+ I1_2_0_1_0_0_0_R0_PLUS I1_2_0_1_1_0_0_R0_MINUS I1_2_0_1_1_0_0_R0_PLUS 
+ I1_2_0_2_0_0_0_R0_MINUS I1_2_0_2_0_0_0_R0_PLUS I1_2_0_2_1_0_0_R0_MINUS 
+ I1_2_0_2_1_0_0_R0_PLUS I1_2_1_0_0_0_0_R0_MINUS I1_2_1_0_0_0_0_R0_PLUS 
+ I1_2_1_0_1_0_0_R0_MINUS I1_2_1_0_1_0_0_R0_PLUS I1_2_1_1_0_0_0_R0_MINUS 
+ I1_2_1_1_0_0_0_R0_PLUS I1_2_1_1_1_0_0_R0_MINUS I1_2_1_1_1_0_0_R0_PLUS 
+ I1_2_1_2_0_0_0_R0_MINUS I1_2_1_2_0_0_0_R0_PLUS I1_2_1_2_1_0_0_R0_MINUS 
+ I1_2_1_2_1_0_0_R0_PLUS I1_2_2_0_0_0_0_R0_MINUS I1_2_2_0_0_0_0_R0_PLUS 
+ I1_2_2_0_1_0_0_R0_MINUS I1_2_2_0_1_0_0_R0_PLUS I1_2_2_1_0_0_0_R0_MINUS 
+ I1_2_2_1_0_0_0_R0_PLUS I1_2_2_1_1_0_0_R0_MINUS I1_2_2_1_1_0_0_R0_PLUS 
+ I1_2_2_2_0_0_0_R0_MINUS I1_2_2_2_0_0_0_R0_PLUS I1_2_2_2_1_0_0_R0_MINUS 
+ I1_2_2_2_1_0_0_R0_PLUS I1_default_MINUS I1_default_PLUS gnd!
*.PININFO I1_0_0_0_0_0_0_R0_MINUS:I I1_0_0_0_0_0_0_R0_PLUS:I 
*.PININFO I1_0_0_0_1_0_0_R0_MINUS:I I1_0_0_0_1_0_0_R0_PLUS:I 
*.PININFO I1_0_0_1_0_0_0_R0_MINUS:I I1_0_0_1_0_0_0_R0_PLUS:I 
*.PININFO I1_0_0_1_1_0_0_R0_MINUS:I I1_0_0_1_1_0_0_R0_PLUS:I 
*.PININFO I1_0_0_2_0_0_0_R0_MINUS:I I1_0_0_2_0_0_0_R0_PLUS:I 
*.PININFO I1_0_0_2_1_0_0_R0_MINUS:I I1_0_0_2_1_0_0_R0_PLUS:I 
*.PININFO I1_0_1_0_0_0_0_R0_MINUS:I I1_0_1_0_0_0_0_R0_PLUS:I 
*.PININFO I1_0_1_0_1_0_0_R0_MINUS:I I1_0_1_0_1_0_0_R0_PLUS:I 
*.PININFO I1_0_1_1_0_0_0_R0_MINUS:I I1_0_1_1_0_0_0_R0_PLUS:I 
*.PININFO I1_0_1_1_1_0_0_R0_MINUS:I I1_0_1_1_1_0_0_R0_PLUS:I 
*.PININFO I1_0_1_2_0_0_0_R0_MINUS:I I1_0_1_2_0_0_0_R0_PLUS:I 
*.PININFO I1_0_1_2_1_0_0_R0_MINUS:I I1_0_1_2_1_0_0_R0_PLUS:I 
*.PININFO I1_0_2_0_0_0_0_R0_MINUS:I I1_0_2_0_0_0_0_R0_PLUS:I 
*.PININFO I1_0_2_0_1_0_0_R0_MINUS:I I1_0_2_0_1_0_0_R0_PLUS:I 
*.PININFO I1_0_2_1_0_0_0_R0_MINUS:I I1_0_2_1_0_0_0_R0_PLUS:I 
*.PININFO I1_0_2_1_1_0_0_R0_MINUS:I I1_0_2_1_1_0_0_R0_PLUS:I 
*.PININFO I1_0_2_2_0_0_0_R0_MINUS:I I1_0_2_2_0_0_0_R0_PLUS:I 
*.PININFO I1_0_2_2_1_0_0_R0_MINUS:I I1_0_2_2_1_0_0_R0_PLUS:I 
*.PININFO I1_1_0_0_0_0_0_R0_MINUS:I I1_1_0_0_0_0_0_R0_PLUS:I 
*.PININFO I1_1_0_0_1_0_0_R0_MINUS:I I1_1_0_0_1_0_0_R0_PLUS:I 
*.PININFO I1_1_0_1_0_0_0_R0_MINUS:I I1_1_0_1_0_0_0_R0_PLUS:I 
*.PININFO I1_1_0_1_1_0_0_R0_MINUS:I I1_1_0_1_1_0_0_R0_PLUS:I 
*.PININFO I1_1_0_2_0_0_0_R0_MINUS:I I1_1_0_2_0_0_0_R0_PLUS:I 
*.PININFO I1_1_0_2_1_0_0_R0_MINUS:I I1_1_0_2_1_0_0_R0_PLUS:I 
*.PININFO I1_1_1_0_0_0_0_R0_MINUS:I I1_1_1_0_0_0_0_R0_PLUS:I 
*.PININFO I1_1_1_0_1_0_0_R0_MINUS:I I1_1_1_0_1_0_0_R0_PLUS:I 
*.PININFO I1_1_1_1_0_0_0_R0_MINUS:I I1_1_1_1_0_0_0_R0_PLUS:I 
*.PININFO I1_1_1_1_1_0_0_R0_MINUS:I I1_1_1_1_1_0_0_R0_PLUS:I 
*.PININFO I1_1_1_2_0_0_0_R0_MINUS:I I1_1_1_2_0_0_0_R0_PLUS:I 
*.PININFO I1_1_1_2_1_0_0_R0_MINUS:I I1_1_1_2_1_0_0_R0_PLUS:I 
*.PININFO I1_1_2_0_0_0_0_R0_MINUS:I I1_1_2_0_0_0_0_R0_PLUS:I 
*.PININFO I1_1_2_0_1_0_0_R0_MINUS:I I1_1_2_0_1_0_0_R0_PLUS:I 
*.PININFO I1_1_2_1_0_0_0_R0_MINUS:I I1_1_2_1_0_0_0_R0_PLUS:I 
*.PININFO I1_1_2_1_1_0_0_R0_MINUS:I I1_1_2_1_1_0_0_R0_PLUS:I 
*.PININFO I1_1_2_2_0_0_0_R0_MINUS:I I1_1_2_2_0_0_0_R0_PLUS:I 
*.PININFO I1_1_2_2_1_0_0_R0_MINUS:I I1_1_2_2_1_0_0_R0_PLUS:I 
*.PININFO I1_2_0_0_0_0_0_R0_MINUS:I I1_2_0_0_0_0_0_R0_PLUS:I 
*.PININFO I1_2_0_0_1_0_0_R0_MINUS:I I1_2_0_0_1_0_0_R0_PLUS:I 
*.PININFO I1_2_0_1_0_0_0_R0_MINUS:I I1_2_0_1_0_0_0_R0_PLUS:I 
*.PININFO I1_2_0_1_1_0_0_R0_MINUS:I I1_2_0_1_1_0_0_R0_PLUS:I 
*.PININFO I1_2_0_2_0_0_0_R0_MINUS:I I1_2_0_2_0_0_0_R0_PLUS:I 
*.PININFO I1_2_0_2_1_0_0_R0_MINUS:I I1_2_0_2_1_0_0_R0_PLUS:I 
*.PININFO I1_2_1_0_0_0_0_R0_MINUS:I I1_2_1_0_0_0_0_R0_PLUS:I 
*.PININFO I1_2_1_0_1_0_0_R0_MINUS:I I1_2_1_0_1_0_0_R0_PLUS:I 
*.PININFO I1_2_1_1_0_0_0_R0_MINUS:I I1_2_1_1_0_0_0_R0_PLUS:I 
*.PININFO I1_2_1_1_1_0_0_R0_MINUS:I I1_2_1_1_1_0_0_R0_PLUS:I 
*.PININFO I1_2_1_2_0_0_0_R0_MINUS:I I1_2_1_2_0_0_0_R0_PLUS:I 
*.PININFO I1_2_1_2_1_0_0_R0_MINUS:I I1_2_1_2_1_0_0_R0_PLUS:I 
*.PININFO I1_2_2_0_0_0_0_R0_MINUS:I I1_2_2_0_0_0_0_R0_PLUS:I 
*.PININFO I1_2_2_0_1_0_0_R0_MINUS:I I1_2_2_0_1_0_0_R0_PLUS:I 
*.PININFO I1_2_2_1_0_0_0_R0_MINUS:I I1_2_2_1_0_0_0_R0_PLUS:I 
*.PININFO I1_2_2_1_1_0_0_R0_MINUS:I I1_2_2_1_1_0_0_R0_PLUS:I 
*.PININFO I1_2_2_2_0_0_0_R0_MINUS:I I1_2_2_2_0_0_0_R0_PLUS:I 
*.PININFO I1_2_2_2_1_0_0_R0_MINUS:I I1_2_2_2_1_0_0_R0_PLUS:I 
*.PININFO I1_default_MINUS:I I1_default_PLUS:I gnd!:I
RI1_2_2_2_1_0_0_R0 I1_2_2_2_1_0_0_R0_PLUS I1_2_2_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=8.0 l=50u w=50u r=6.53672 par=8.0 s=1
RI1_2_2_2_0_0_0_R0 I1_2_2_2_0_0_0_R0_PLUS I1_2_2_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=50u w=50u r=6.53672 par=1.0 s=8
RI1_2_2_1_1_0_0_R0 I1_2_2_1_1_0_0_R0_PLUS I1_2_2_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=3.0 l=50u w=50u r=6.53672 par=3.0 s=1
RI1_2_2_1_0_0_0_R0 I1_2_2_1_0_0_0_R0_PLUS I1_2_2_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=50u w=50u r=6.53672 par=1.0 s=3
RI1_2_2_0_1_0_0_R0 I1_2_2_0_1_0_0_R0_PLUS I1_2_2_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=50u w=50u r=6.53672 par=1.0 s=1
RI1_2_2_0_0_0_0_R0 I1_2_2_0_0_0_0_R0_PLUS I1_2_2_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=50u w=50u r=6.53672 par=1.0 s=1
RI1_2_1_2_1_0_0_R0 I1_2_1_2_1_0_0_R0_PLUS I1_2_1_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=8.0 l=2.6u w=50u r=567.308m par=8.0 s=1
RI1_2_1_2_0_0_0_R0 I1_2_1_2_0_0_0_R0_PLUS I1_2_1_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=2.6u w=50u r=567.308m par=1.0 s=8
RI1_2_1_1_1_0_0_R0 I1_2_1_1_1_0_0_R0_PLUS I1_2_1_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=3.0 l=2.6u w=50u r=567.308m par=3.0 s=1
RI1_2_1_1_0_0_0_R0 I1_2_1_1_0_0_0_R0_PLUS I1_2_1_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=2.6u w=50u r=567.308m par=1.0 s=3
RI1_2_1_0_1_0_0_R0 I1_2_1_0_1_0_0_R0_PLUS I1_2_1_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=2.6u w=50u r=567.308m par=1.0 s=1
RI1_2_1_0_0_0_0_R0 I1_2_1_0_0_0_0_R0_PLUS I1_2_1_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=2.6u w=50u r=567.308m par=1.0 s=1
RI1_2_0_2_1_0_0_R0 I1_2_0_2_1_0_0_R0_PLUS I1_2_0_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=8.0 l=840n w=50u r=345.658m par=8.0 s=1
RI1_2_0_2_0_0_0_R0 I1_2_0_2_0_0_0_R0_PLUS I1_2_0_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=840n w=50u r=345.658m par=1.0 s=8
RI1_2_0_1_1_0_0_R0 I1_2_0_1_1_0_0_R0_PLUS I1_2_0_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=3.0 l=840n w=50u r=345.658m par=3.0 s=1
RI1_2_0_1_0_0_0_R0 I1_2_0_1_0_0_0_R0_PLUS I1_2_0_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=840n w=50u r=345.658m par=1.0 s=3
RI1_2_0_0_1_0_0_R0 I1_2_0_0_1_0_0_R0_PLUS I1_2_0_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=840n w=50u r=345.658m par=1.0 s=1
RI1_2_0_0_0_0_0_R0 I1_2_0_0_0_0_0_R0_PLUS I1_2_0_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=840n w=50u r=345.658m par=1.0 s=1
RI1_1_2_2_1_0_0_R0 I1_1_2_2_1_0_0_R0_PLUS I1_1_2_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=8.0 l=50u w=1.57u r=205.015 par=8.0 s=1
RI1_1_2_2_0_0_0_R0 I1_1_2_2_0_0_0_R0_PLUS I1_1_2_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=50u w=1.57u r=205.015 par=1.0 s=8
RI1_1_2_1_1_0_0_R0 I1_1_2_1_1_0_0_R0_PLUS I1_1_2_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=3.0 l=50u w=1.57u r=205.015 par=3.0 s=1
RI1_1_2_1_0_0_0_R0 I1_1_2_1_0_0_0_R0_PLUS I1_1_2_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=50u w=1.57u r=205.015 par=1.0 s=3
RI1_1_2_0_1_0_0_R0 I1_1_2_0_1_0_0_R0_PLUS I1_1_2_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=50u w=1.57u r=205.015 par=1.0 s=1
RI1_1_2_0_0_0_0_R0 I1_1_2_0_0_0_0_R0_PLUS I1_1_2_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=50u w=1.57u r=205.015 par=1.0 s=1
RI1_1_1_2_1_0_0_R0 I1_1_1_2_1_0_0_R0_PLUS I1_1_1_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=8.0 l=2.6u w=1.57u r=17.7928 par=8.0 s=1
RI1_1_1_2_0_0_0_R0 I1_1_1_2_0_0_0_R0_PLUS I1_1_1_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=2.6u w=1.57u r=17.7928 par=1.0 s=8
RI1_1_1_1_1_0_0_R0 I1_1_1_1_1_0_0_R0_PLUS I1_1_1_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=3.0 l=2.6u w=1.57u r=17.7928 par=3.0 s=1
RI1_1_1_1_0_0_0_R0 I1_1_1_1_0_0_0_R0_PLUS I1_1_1_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=2.6u w=1.57u r=17.7928 par=1.0 s=3
RI1_1_1_0_1_0_0_R0 I1_1_1_0_1_0_0_R0_PLUS I1_1_1_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=2.6u w=1.57u r=17.7928 par=1.0 s=1
RI1_1_1_0_0_0_0_R0 I1_1_1_0_0_0_0_R0_PLUS I1_1_1_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=2.6u w=1.57u r=17.7928 par=1.0 s=1
RI1_1_0_2_1_0_0_R0 I1_1_0_2_1_0_0_R0_PLUS I1_1_0_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=8.0 l=840n w=1.57u r=10.8411 par=8.0 s=1
RI1_1_0_2_0_0_0_R0 I1_1_0_2_0_0_0_R0_PLUS I1_1_0_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=840n w=1.57u r=10.8411 par=1.0 s=8
RI1_1_0_1_1_0_0_R0 I1_1_0_1_1_0_0_R0_PLUS I1_1_0_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=3.0 l=840n w=1.57u r=10.8411 par=3.0 s=1
RI1_1_0_1_0_0_0_R0 I1_1_0_1_0_0_0_R0_PLUS I1_1_0_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=840n w=1.57u r=10.8411 par=1.0 s=3
RI1_1_0_0_1_0_0_R0 I1_1_0_0_1_0_0_R0_PLUS I1_1_0_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=840n w=1.57u r=10.8411 par=1.0 s=1
RI1_1_0_0_0_0_0_R0 I1_1_0_0_0_0_0_R0_PLUS I1_1_0_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=840n w=1.57u r=10.8411 par=1.0 s=1
RI1_0_2_2_1_0_0_R0 I1_0_2_2_1_0_0_R0_PLUS I1_0_2_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=8.0 l=50u w=420n r=734.83 par=8.0 s=1
RI1_0_2_2_0_0_0_R0 I1_0_2_2_0_0_0_R0_PLUS I1_0_2_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=50u w=420n r=734.83 par=1.0 s=8
RI1_0_2_1_1_0_0_R0 I1_0_2_1_1_0_0_R0_PLUS I1_0_2_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=3.0 l=50u w=420n r=734.83 par=3.0 s=1
RI1_0_2_1_0_0_0_R0 I1_0_2_1_0_0_0_R0_PLUS I1_0_2_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=50u w=420n r=734.83 par=1.0 s=3
RI1_0_2_0_1_0_0_R0 I1_0_2_0_1_0_0_R0_PLUS I1_0_2_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=50u w=420n r=734.83 par=1.0 s=1
RI1_0_2_0_0_0_0_R0 I1_0_2_0_0_0_0_R0_PLUS I1_0_2_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=50u w=420n r=734.83 par=1.0 s=1
RI1_0_1_2_1_0_0_R0 I1_0_1_2_1_0_0_R0_PLUS I1_0_1_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=8.0 l=2.6u w=420n r=63.7743 par=8.0 s=1
RI1_0_1_2_0_0_0_R0 I1_0_1_2_0_0_0_R0_PLUS I1_0_1_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=2.6u w=420n r=63.7743 par=1.0 s=8
RI1_0_1_1_1_0_0_R0 I1_0_1_1_1_0_0_R0_PLUS I1_0_1_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=3.0 l=2.6u w=420n r=63.7743 par=3.0 s=1
RI1_0_1_1_0_0_0_R0 I1_0_1_1_0_0_0_R0_PLUS I1_0_1_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=2.6u w=420n r=63.7743 par=1.0 s=3
RI1_0_1_0_1_0_0_R0 I1_0_1_0_1_0_0_R0_PLUS I1_0_1_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=2.6u w=420n r=63.7743 par=1.0 s=1
RI1_0_1_0_0_0_0_R0 I1_0_1_0_0_0_0_R0_PLUS I1_0_1_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=2.6u w=420n r=63.7743 par=1.0 s=1
RI1_0_0_2_1_0_0_R0 I1_0_0_2_1_0_0_R0_PLUS I1_0_0_2_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=8.0 l=840n w=420n r=38.8574 par=8.0 s=1
RI1_0_0_2_0_0_0_R0 I1_0_0_2_0_0_0_R0_PLUS I1_0_0_2_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=840n w=420n r=38.8574 par=1.0 s=8
RI1_0_0_1_1_0_0_R0 I1_0_0_1_1_0_0_R0_PLUS I1_0_0_1_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=3.0 l=840n w=420n r=38.8574 par=3.0 s=1
RI1_0_0_1_0_0_0_R0 I1_0_0_1_0_0_0_R0_PLUS I1_0_0_1_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=840n w=420n r=38.8574 par=1.0 s=3
RI1_0_0_0_1_0_0_R0 I1_0_0_0_1_0_0_R0_PLUS I1_0_0_0_1_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=840n w=420n r=38.8574 par=1.0 s=1
RI1_0_0_0_0_0_0_R0 I1_0_0_0_0_0_0_R0_PLUS I1_0_0_0_0_0_0_R0_MINUS $SUB=gnd! 
+ $[nplus_s_dw] m=1.0 l=840n w=420n r=38.8574 par=1.0 s=1
RI1_default I1_default_PLUS I1_default_MINUS $SUB=gnd! $[nplus_s_dw] m=1.0 
+ l=840.00n w=420.00n r=38.8574 par=1.0 s=1
.ENDS

