.SUBCKT gf180mcu_fd_io__brk5 VSS
.ENDS
