***************************
** pfet_03v3_t_id
***************************
* Copyright 2022 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
Vds D_tn 0 dc -3.3
Vgs G_tn 0 -3.3

.temp {{temp}}
 
xmn1 D_tn G_tn 0 0 {{device}} W = {{width}}u L = {{length}}u

**** begin architecture code

.control
set filetype=ascii
set wr_singlescale
set wr_vecnames
dc Vds {{vds}} Vgs {{vgs}}

wrdata mos_iv_regr/{{device}}/{{device}}_netlists_Id/T{{temp}}_simulated_W{{width}}_L{{length}}.csv i(Vds) v(G_tn) v(D_tn) 
.endc

** library calling

.include "../../../design.ngspice"
.lib "../../../sm141064.ngspice" typical

**** end architecture code

.end
