*****************
** main netlist
*****************

Vcp c 0 dc 3
Vbp b 0 dc 1.2

xq1 c b 0 0 {{device}}


*****************
** Analysis
*****************
.control

.DC Vbp 0.2 1.2 0.01 Vcp 1 3 1
.STEP TEMP {{temp}} -60 200

.print DC FORMAT=CSV file=bjt_beta_reg/npn/simulated_Ic/t{{temp}}_simulated_{{device}}.csv {-I(Vcp)} v(b) v(c)



.include "../../../design.xyce"
.lib "../../../sm141064.xyce" bjt_typical

.end
