***************************
** nfet_03v3_t_id
***************************
* Copyright 2022 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

** library calling

.include "../../../design.ngspice"
.lib "../../../sm141064.ngspice" typical



** Circuit Description **
* power supply
vds D_tn 0 dc=0
vgs G_tn 0 dc=3.3
vbs S_tn 0 dc=0

.temp 25
.options tnom=25


* circuit
mn 0 G_tn 0 S_tn {{device}} W = {{width}}u L = {{length}}u nf={{nf}} ad={{AD}}u pd={{PD}}u as={{AS}}u ps={{PS}}u

.control
set filetype=ascii
set wr_singlescale
set wr_vecnames

compose  vbs_vector   start={{vbs1}}          stop={{vbs2}}          step={{vbs3}}

set appendwrite

foreach t 25

    let vbs_counter = 0
    while vbs_counter < length(vbs_vector)
        option TEMP=25
        alter vbs = vbs_vector[vbs_counter]

        save  @mn[vs] @mn[vgs] @mn[id] @mn[cgb]
        *******************
        ** simulation part
        *******************
        DC vgs {{vgs}}
    
        * ** parameters calculation
	
	let Cap = -{@mn[cgb]*1e15}
        let Vg = -1*@mn[vbs]
        
        wrdata mos_cv_regr/{{device}}/{{device}}_netlists_Cgc/simulated_W{{width}}_L{{length}}.csv Cap Vg
        
        reset
        let vbs_counter = vbs_counter + 1
    end
end
.endc
.end
