*Xyce Common Source Circuit
** library calling


*****************
** main netlist
*****************
Vn n 0 dc 1

*r1 n p 1MEG
xrn n 0 0 ppolyf_s L=50u W=150u
* PJ=40u

* .print dc Rs=par('(1M*V(p)/(V(n)-V(p)))/100u*100u')

*****************
** Analysis
*****************
.OP
* .DC Vn 1 1 0.1
* .print DC FORMAT=CSV file=result.csv {(1MEG*V(p)/(V(n)-V(p)))/50u*150u}
.print DC FORMAT=CSV file=result.csv {(V(n)*150u)/(-I(Vn)*50u)}


.include "../../../../design.xyce"
.lib "../../../../sm141064.xyce" res_typical

.end