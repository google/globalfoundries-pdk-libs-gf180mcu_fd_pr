*Xyce Common Source Circuit
** library calling



*****************
** main netlist
*****************
Vds D_tn 0 dc 3.3
Vgs G_tn 0 dc 3.3


xmn1 D_tn G_tn 0 0 {{device}} W={{width}}u L={{length}}u ad={{AD}}u pd={{PD}}u as={{AS}}u ps={{PS}}u

*****************
** Analysis
*****************
.DC Vds {{vds}} Vgs {{vgs}}
.STEP TEMP {{temp}} -60 200
.print DC FORMAT=CSV file=mos_iv_reg/{{device}}/{{device}}_netlists_Id/t{{temp}}_simulated_W{{width}}_L{{length}}.csv {-I(Vds)} v(D_tn) v(G_tn)

.include "../../../../../../design.xyce"
.lib "../../../../../../sm141064.xyce" typical

.end
