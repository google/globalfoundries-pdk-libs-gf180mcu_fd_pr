*Xyce Common Source Circuit
** library calling


*****************
** main netlist
*****************
Vds D_tn 0 dc 0.05
Vgs G_tn 0 dc 3.3
Vbs B_tn 0 dc 0

xmn1 D_tn G_tn 0 B_tn {{device}} W={{width}}u L={{length}}u ad={{AD}}u pd={{PD}}u as={{AS}}u ps={{PS}}u


*****************
** Analysis
*****************
.dc Vgs {{vgs}} Vbs {{vbs}}
.STEP TEMP {{temp}} -60 200
.print DC FORMAT=CSV file=mos_iv_reg/{{device}}/{{device}}_netlists_Id/t{{temp}}_simulated_W{{width}}_L{{length}}.csv {-I(Vds)} v(G_tn) v(B_tn)

.include "../../../../../../design.xyce"
.lib "../../../../../../sm141064.xyce" typical

.end
