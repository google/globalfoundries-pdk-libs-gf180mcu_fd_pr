***************************
** CV netlist generation **
***************************
* Copyright 2022 Efabless Corporation
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
Vn n 0 dc 1


.temp {{temp}}
.options tnom={{temp}}
      

dn n 0 {{device}} AREA = {{area}}p PJ = {{pj}}u 

.control
set filetype=ascii

let vn_min  = 0
let vn_step = -0.2
let vn_max  = -3.2

option TEMP={{temp}}

save   @dn[cd]
*******************
** simulation part
*******************
DC Vn $&vn_min $&vn_max $&vn_step

* ** parameters calculation

print  @dn[cd]*1000000000000000
    
wrdata diode_regr/{{device}}/{{device}}_netlists_cv/simulated_W{{width}}_L{{length}}_t{{temp}}_{{corner}}.csv  @dn[cd]*1000000000000000


.endc

** library calling

.include "../../../design.ngspice"
.lib "../../../sm141064.ngspice" diode_{{corner}}


.end
